------ shifter_map1

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

ENTITY S_MAP1 IS
GENERIC(
		n : INTEGER := 16;
		addr_col  : integer := 10; -- required bits to store 16 elements
		col : integer := 1023; --- = H
        addr_row  : integer := 4; -- required bits to store 16 elements
		row : integer :=12 -- = n
        );
PORT ( 
      clk, rst, run: in std_logic;
      reg_out : out std_logic;
      din :in std_logic_vector(15 downto 0);
      df , do , dc ,di : out std_logic_vector (31 downto 0)
	   );
END S_MAP1;	  


ARCHITECTURE behavioral OF S_MAP1 IS

component ROM is
    generic(
        addr_col  : integer := 10; -- required bits to store 16 elements
		col : integer := 1023;
        addr_row  : integer := 4; -- required bits to store 16 elements
		row : integer :=12
        );
	port(
		addr_c : in std_logic_vector(addr_col downto 0);
		addr_r : in std_logic_vector(addr_row downto 0);
		data : out std_logic_vector(19 downto 0)
	);
end component;

component single_port_RAM is
  generic ( n : integer := 15;
			addr_width : integer := 4 ;
			row : integer := 4 
			);
  port(
    clk: in std_logic;
    we : in std_logic;
    addr : in std_logic_vector(addr_row downto 0);
    din : in std_logic_vector(n downto 0);
    dout : out std_logic_vector(n downto 0)
    );
end component;

component map_shifter_controller IS
  generic ( 
		n : INTEGER := 16;
		addr_col  : INTEGER := 8; -- required bits to store 16 elements
		col : INTEGER := 350;
        addr_row  : INTEGER := 4; -- required bits to store 16 elements
		row : INTEGER :=8 
		);
  PORT ( 
      clk, rst, run : in STD_LOGIC;
      add_reg, out_reg, we_input_reg :out STD_LOGIC ;
	  add_row : out STD_LOGIC_VECTOR (addr_row downto 0);
	  add_col : out STD_LOGIC_VECTOR (addr_col downto 0));  
END component;

component mul IS
  PORT ( 
      s1, s2, s3, s4 :in STD_LOGIC;
      load1, load2, load3, load4 : in STD_LOGIC_VECTOR(3 downto 0);
      din : in STD_LOGIC_VECTOR(15 downto 0);
	  dout1, dout2, dout3, dout4 : out STD_LOGIC_VECTOR(15 downto 0));
END component;    
    
component cla_4 IS
	PORT ( 
		  clk, rst, add_reg, out_reg: in std_logic;
		  mulx1, mulx2, mulx3, mulx4 : in std_logic_vector (15 downto 0);
		  df , do , dc ,di : out std_logic_vector (31 downto 0)
		   );
END component;

signal addr_r :  STD_LOGIC_VECTOR (addr_row downto 0);
signal addr_c : STD_LOGIC_VECTOR (addr_col downto 0);
signal add_reg, out_reg , we: std_logic;
signal wf,wo, wi , wc :std_logic_vector(3 downto 0);
signal sx1, sx2, sx3, sx4 :std_logic;
signal mulx1, mulx2, mulx3, mulx4, dout :std_logic_vector(15 downto 0);
signal data : std_logic_vector(19 downto 0);
signal dfm , dom , dcm ,dim : std_logic_vector (31 downto 0);

BEGIN

MAP1_ROM : ROM 
    generic MAP(
        addr_col ,
		col ,
        addr_row ,
		row )
	port MAP(
		addr_c ,
		addr_r ,
		data );
	
INPUT_RAM : single_port_RAM
  generic MAP( 
			15,
			addr_row ,
			row
			)
  port MAP(
    clk, we, addr_r , din, dout   );

control : map_shifter_controller
  generic map (n ,addr_col ,col ,addr_row  ,row ) 
  port map(
      clk, rst, run ,
      add_reg, out_reg,we,
	  addr_r, addr_c
	   );
	  
mull_shift : mul 
  port map(
      sx1, sx2, sx3, sx4 ,
      wf,wo, wi , wc ,
      dout,
	  mulx1, mulx2, mulx3, mulx4 );
	  
adding_map : cla_4 
	PORT map( 
		  clk, rst, add_reg, out_reg,
		  mulx1, mulx2, mulx3, mulx4,
		  dfm , dom , dcm ,dim
		   );
	df <= dfm;
	do <= dom;
	dc <= dcm;
	di <= dim;
	sx1 <=data(4);
    sx2 <=data(9);
    sx3 <=data(14);
    sx4 <=data(19);
    wf <=data(3 downto 0);
    wo <=data(8 downto 5);
    wi <=data(13 downto 10);
    wc <=data(18 downto 15);
	reg_out <= out_reg;
END behavioral;	 
-----------------------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

ENTITY cla_4 IS
	PORT ( 
		  clk, rst, add_reg, out_reg: in std_logic;
		  mulx1, mulx2, mulx3, mulx4 : in std_logic_vector (15 downto 0);
		  df , do , dc ,di : out std_logic_vector (31 downto 0)
		   );
END cla_4;	  


ARCHITECTURE behavioral OF cla_4 IS
    
component add_cla IS
  PORT ( 
      clk, rst,  add_reg, out_reg: in STD_LOGIC;
      din1 : in STD_LOGIC_VECTOR(15 downto 0);
	  dout : out STD_LOGIC_VECTOR(31 downto 0));
END component;

BEGIN

addf : add_cla 
  port map(
      clk, rst, add_reg, out_reg,
      mulx1, 
	  df );
addc : add_cla 
  port map(
      clk, rst, add_reg, out_reg,
      mulx2,
	  dc );
addi : add_cla 
  port map(
      clk, rst, add_reg, out_reg,
      mulx3, 
	  di );
addo : add_cla 
  port map(
      clk, rst, add_reg, out_reg,
      mulx4,
	  do );

END behavioral;	 
-----------------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

ENTITY mul IS
PORT (s1, s2, s3, s4 :in STD_LOGIC;
      load1, load2, load3, load4 : in STD_LOGIC_VECTOR(3 downto 0);
      din : in STD_LOGIC_VECTOR(15 downto 0);
	  dout1, dout2, dout3, dout4 : out STD_LOGIC_VECTOR(15 downto 0));
END mul;	  

ARCHITECTURE behavioral OF mul Is
signal l1 , l2 , l3 , l4 : integer ;
BEGIN
		--l1 <=16 - to_integer(unsigned(load1));
		--l2 <=16 - to_integer(unsigned(load2));
		--l3 <=16 - to_integer(unsigned(load3));
		--l4 <=16 - to_integer(unsigned(load4));
		dout1(14 downto 0)<= std_logic_vector( shift_right( unsigned(din(14 downto 0)),to_integer(unsigned(load1))));
		dout2(14 downto 0)<= std_logic_vector( shift_right( unsigned(din(14 downto 0)),to_integer(unsigned(load2))));
		dout3(14 downto 0)<= std_logic_vector( shift_right( unsigned(din(14 downto 0)),to_integer(unsigned(load3))));
		dout4(14 downto 0)<= std_logic_vector( shift_right( unsigned(din(14 downto 0)),to_integer(unsigned(load4))));
        dout1(15) <= s1 xor din(15);
        dout2(15) <= s2 xor din(15);
        dout3(15) <= s3 xor din(15);
        dout4(15) <= s4 xor din(15);
END behavioral;	 

------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;

ENTITY map_shifter_controller IS
generic(
		n : INTEGER := 16;
		addr_col  : INTEGER := 4; -- required bits to store 16 elements
		col : INTEGER := 16;
        addr_row  : INTEGER := 4; -- required bits to store 16 elements
		row : INTEGER :=16 ); -- = n
PORT ( 
	clk, rst, run : in STD_LOGIC;
	add_reg, out_reg, we_input_reg :out STD_LOGIC ;
	add_row : out STD_LOGIC_VECTOR (addr_row downto 0);
	add_col : out STD_LOGIC_VECTOR (addr_col downto 0)
  );       
END map_shifter_controller;	  

ARCHITECTURE contr OF map_shifter_controller Is

component counter IS
	generic ( n : INTEGER := 8);
	PORT ( 
		  clk, rst,  en: in STD_LOGIC;
		  dout : out STD_LOGIC_VECTOR(n downto 0));
END component;

  signal add_row_i , r_i : STD_LOGIC_VECTOR (addr_row downto 0);
  signal add_col_i , c_i: STD_LOGIC_VECTOR (addr_col downto 0);
  TYPE mini_state IS  (init, wait_s,rst_mull_count1,rst_mull_count2,  mull,  end_reg,  end_reg_f); -- add_pause,  
  SIGNAL ns,  ps : mini_state;
  SIGNAL count_r , rst_count_r, count_c , rst_count_c : STD_LOGIC;
  
BEGIN 
-- c <= STD_LOGIC_VECTOR(to_UNSIGNED(n , 4));
PROCESS(clk) BEGIN 
  IF rising_edge(clk) then
    IF (rst ='1')then
      ps <= init; 
    ELSe  
      ps <= ns;  
    END IF;
  END IF;
END PROCESS;

PROCESS ( ps,  run,  add_row_i, add_col_i )
  BEGIN 
    add_reg <= '0';
    out_reg <= '0';
	count_r <= '0';
	count_c <= '0';
	rst_count_c <= '0';
	rst_count_r <= '0';
	we_input_reg <= '0';
  CASE (ps) IS 
    WHEN init => 
		rst_count_c <= '1';
		rst_count_r <= '1';
		IF ( run = '1') then
			ns <= wait_s;
        ELSe
			ns <= init;
        END IF;
	WHEN wait_s => 
		we_input_reg <= '1';
		count_r <= '1';
		IF ( add_row_i = r_i) then 
			ns <= rst_mull_count1;
		ELSe 
			ns <= wait_s;
		END IF;
	when rst_mull_count1 =>
		rst_count_r <= '1';
			ns <= mull;
    WHEN mull =>
		count_r <= '1';
		add_reg <= '1';
		IF ( add_row_i = r_i) then 
			ns <= end_reg;
		ELSe 
			ns <= mull;
		END IF;
    WHEN end_reg =>
		count_c <= '1';
		out_reg <= '1';
		rst_count_r <= '1';
		IF ( add_col_i = c_i) then 
			ns <= end_reg_f;
		ELSe 
			ns <= mull;
		END IF;
	WHEN end_reg_f =>
		rst_count_r <= '1';
		rst_count_c <= '1';
		IF ( run = '1') then
			ns <= wait_s;
        ELSe
			ns <= init;
        END IF;
    WHEN OTHERS =>
			ns <= init;
   END CASE;
END PROCESS;
 
c_count : counter 
	generic map(addr_col)
	PORT map( 
		  clk, rst_count_c,  count_c ,add_col_i);
r_count : counter 
	generic map(addr_row)
	PORT map( 
		  clk, rst_count_r, count_r , add_row_i);
	r_i <= STD_LOGIC_VECTOR(to_UNSIGNED((row -1), addr_row+1));
	c_i <= STD_LOGIC_VECTOR(to_UNSIGNED((col -1), addr_col+1));
	add_col <= add_col_i;
	add_row <= add_row_i;
		  
END contr;	 
------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY counter IS
generic ( n : integer := 8);
PORT ( 
      clk, rst,  en: in STD_LOGIC;
	  dout : out STD_LOGIC_VECTOR(n downto 0));
END counter;	  

ARCHITECTURE behavioral OF counter IS
signal i : std_logic_vector(n downto 0);
begin
PROCESS (clk)
	   BEGIN 
		 IF rising_edge (clk ) then 
		     IF ( rst = '1') then 
			 	i <= (others => '0'); 
		     ELSIF ( en = '1')then
		        i <= STD_LOGIC_VECTOR(UNSIGNED(i)+ 1);
		     END IF;
	     END IF;
END PROCESS;
dout <= i ; 
end behavioral;
  
------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY add_cla IS
PORT ( 
      clk, rst,  add_reg, out_reg: in STD_LOGIC;
      din1 : in STD_LOGIC_VECTOR(15 downto 0);
	  dout : out STD_LOGIC_VECTOR(31 downto 0));
END add_cla;	  

ARCHITECTURE behavioral OF add_cla IS
  
component  cla_add_16_32 IS
PORT (  din1, din2 : in STD_LOGIC_VECTOR(31 downto 0);
	    dout : out STD_LOGIC_VECTOR(31 downto 0));
END component;


signal outm1, d, d_reg2, outreg : std_logic_vector(31 downto 0);

BEGIN

 d <= din1(15)& "0000000000000000"& din1(14 downto 0);

 PROCESS(clk)
	 BEGIN 
	   IF rising_edge(clk )THEN
	     IF (rst ='1') THEN
			d_reg2 <= (OTHERS => '0');
			outreg <= (OTHERS => '0');
		 ELSIF (add_reg = '1')THEN
			d_reg2 <= outm1;
			outreg <= outreg;
		 ELSIF (out_reg ='1') THEN
			outreg <= d_reg2;
			d_reg2 <= (OTHERS =>'0');
		 ELSE
			d_reg2 <= d_reg2;
			outreg <= outreg;
		 END IF; 
	   END IF;
	END PROCESS;  

add1 : cla_add_16_32 
      port map ( d , d_reg2 , outm1);  

dout <= outreg; 

END behavioral;	
---------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use IEEE.numeric_std.all; 

ENTITY cla_add_16_32 IS
PORT (din1, din2 : in STD_LOGIC_VECTOR(31 downto 0);
	    dout : out STD_LOGIC_VECTOR(31 downto 0));
END cla_add_16_32;	  

ARCHITECTURE behavioral OF cla_add_16_32 IS

signal out1, out2, d : std_logic_vector(31 downto 0);
signal en , se11, sel2, sign : std_logic;
--signal val : std_logic_vector(31 downto 0):= (others =>'0');
signal do : std_logic_vector(31 downto 0);


component twoscompliment IS
generic ( n : integer := 31);
PORT (en : in std_logic;
      din : in STD_LOGIC_VECTOR(n downto 0);
	    dout : out STD_LOGIC_VECTOR(n downto 0));
END component;

component mux_2 is
  generic (
		n : integer := 31
		);
  port (
        sel : in std_logic;
        a , b : in STD_LOGIC_VECTOR (n DOWNTO 0);
        c :out STD_LOGIC_VECTOR(n DOWNTO 0) 
         );
end component;

component cla_16_32 IS
PORT ( din1, din2 : in STD_LOGIC_VECTOR(31 downto 0);
       dout : out STD_LOGIC_VECTOR(31 downto 0));
END component;

BEGIN
    
process(din1,din2)
 begin
  
    if ( din1(31) = din2(31) ) then
       en <= '0';
       se11 <= '0'; -- din1
       sel2 <= '1'; -- din2
       --sign <= din1(31);
    ELSif (din1(30 downto 0) > din2(30 downto 0)) then
       en <= '1';
       se11 <= '0'; -- din1
       sel2 <= '1'; -- din2
       --sign <= din1(31);
    else
       en <= '1';
       se11 <= '1'; -- din1
       sel2 <= '0'; -- din2
      -- sign <= din2(31);
    end if;
    
 end process;
 
 comp : twoscompliment 
	generic map (31)
    PORT MAP(en ,
      out2 ,
	    d);
	    
  mux0 :mux_2 
  generic map (31)
  port map(
        se11 ,
        din1 , din2,
        out1
         );
  mux1 :mux_2 
  generic map (31)
  port map(
        sel2 ,
        din1 , din2,
        out2
         );      
  adding : cla_16_32
  PORT MAP ( out1, d , do);
  
  dout  <= do(31 downto 0);
  
END behavioral;
--------------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY add IS
PORT ( 
      clk, rst,  add_reg, out_reg: in STD_LOGIC;
      din1 : in STD_LOGIC_VECTOR(15 downto 0);
	  dout : out STD_LOGIC_VECTOR(31 downto 0));
END add;	  

ARCHITECTURE behavioral OF add IS
  
component  cla_add_16_32 IS
PORT (  din1, din2 : in STD_LOGIC_VECTOR(31 downto 0);
	    dout : out STD_LOGIC_VECTOR(31 downto 0));
END component;


signal outm1, d, d_reg2, outreg : std_logic_vector(31 downto 0);

BEGIN

 d <= din1(15)& "0000000000000000"& din1(14 downto 0);

 PROCESS(clk)
	 BEGIN 
	   IF rising_edge(clk )THEN
	     IF (rst ='1') THEN
			d_reg2 <= (OTHERS => '0');
			outreg <= (OTHERS => '0');
		 ELSIF (add_reg = '1')THEN
			d_reg2 <= outm1;
			outreg <= outreg;
		 ELSIF (out_reg ='1') THEN
			outreg <= d_reg2;
			d_reg2 <= (OTHERS =>'0');
		 ELSE
			d_reg2 <= d_reg2;
			outreg <= outreg;
		 END IF; 
	   END IF;
	END PROCESS;  

add1 : cla_add_16_32 
      port map ( d , d_reg2 , outm1);  

dout <= outreg; 

END behavioral;	
------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY CLG_16 IS
PORT ( p,g,a: in STD_LOGIC_VECTOR(15 downto 0);
      c0 : in std_logic;
       c : out STD_LOGIC_VECTOR(15 downto 0));
END CLG_16;	  

ARCHITECTURE behavioral OF CLG_16 IS
signal x0, x1, x2, x3, x4 , x5, x6, x7, x8,x9,x10, x11, x12, x13, x14 , x15, x16 : std_logic;
signal y0, y1, y2, y3, y4 , y5, y6, y7, y8,y9,y10, y11, y12, y13, y14 , y15 : std_logic;
signal z0, z1, z2, z3, z4 , z5, z6, z7, z8,z9,z10, z11, z12, z13, z14 , z15 : std_logic;
BEGIN
  x0 <= a(0) and c0;
  x1 <= a(1) and x0;
  x2 <= a(2) and x1;
  x3 <= a(3) and x2;
  x4 <= a(4) and x3;
  x5 <= a(5) and x4;
  x6 <= a(6) and x5;
  x7 <= a(7) and x6;
  x8 <= a(8) and x7;
  x9 <= a(9) and x8;
  x10 <= a(10) and x9;
  x11 <= a(11) and x10;
  x12 <= a(12) and x11;
  x13 <= a(13) and x12;
  x14 <= a(14) and x13;
  x15 <= a(15) and x14;
  y0 <= a(1) and g(0);
  y1 <= a(2) and y0;
  y2 <= a(3) and y1;
  y3 <= a(4) and y2;
  y4 <= a(5) and y3;
  y5 <= a(6) and y4;
  y6 <= a(7) and y5;
  y7 <= a(8) and y6;
  y8 <= a(9) and y7;
  y9 <= a(10) and y8;
  y10 <= a(11) and y9;
  y11 <= a(12) and y10;
  y12 <= a(13) and y11;
  y13 <= a(14) and y12;
  y14 <= a(15) and y13;

 c(0) <= g(0) or x0;
   c(1) <= g(1) or y0 or x1;
   c(2) <= g(2) or (a(2) and g(1)) or y1 or x2;
   c(3) <= g(3) or (a(3) and g(2)) or (a(3) and a(2) and g(1)) or y2 or x3;
   c(4) <= g(4) or (a(4) and g(3)) or (a(4) and a(3) and g(2)) or (a(4) and a(3) and a(2) and g(1)) or y3 or x4;
   c(5) <= g(5) or (a(5) and g(4)) or (a(5) and a(4) and g(3)) or (a(5) and a(4) and a(3) and g(2)) or y4 or x5;
   c(6) <= g(6) or (a(6) and g(5)) or (a(6) and a(5) and g(4)) or (a(6) and a(5) and a(4) and g(3)) or (a(6) and a(5) and a(4) and a(3) and g(2)) or y5 or x6;
    c(7) <= g(7) or (a(7) and g(6)) or (a(7) and a(6) and g(5)) or (a(7) and a(6) and a(5) and g(4)) or (a(7) and a(6) and a(5) and a(4) and g(3)) or (a(7) and a(6) and a(5) and a(4) and 
                a(3) and g(2)) or (a(7) and a(6) and a(5) and a(4) and a(3) and a(2)  and g(1)) or y6 or x7;
    c(8) <= g(8) or (a(8) and g(7)) or (a(8) and a(7) and g(6)) or (a(8) and a(7) and a(6) and g(5)) or (a(8) and a(7) and a(6) and a(5)  and g(4)) or (a(8) and a(7) and a(6) and a(5) and a(4)  
                 and g(3)) or (a(8) and a(7) and a(6) and a(5) and a(4) and a(3)   and g(2)) or (a(8) and a(7) and a(6) and a(5) and a(4) and a(3) and a(2)   and g(1)) or y7 or x8;
     c(9) <= g(9) or (a(9) and g(8)) or (a(9) and a(8) and g(7)) or (a(9) and a(8) and a(7)  and g(6)) or (a(9) and a(8) and a(7) and a(6)  and g(5)) or (a(9) and a(8) and a(7) and a(6) and a(5)   
                 and g(4)) or (a(9) and a(8) and a(7) and a(6) and a(5) and a(4)  and g(3)) or (a(9) and a(8) and a(7) and a(6) and a(5) and a(4) and a(3)  and g(2)) or (a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y8 or  x9;
     c(10) <= g(10) or (a(10) and g(9)) or (a(10) and a(9) and g(8)) or (a(10) and a(9) and a(8)  and g(7)) or (a(10) and a(9) and a(8) and a(7)  and g(6)) or (a(10) and a(9) and a(8) and a(7) and a(6)   
                 and g(5)) or (a(10) and a(9) and a(8) and a(7) and a(6) and a(5) and g(4)) or (a(10) and a(9) and a(8) and a(7) and a(6) and a(5) and a(4) and g(3)) or (a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and g(2)) or (a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y9 or x10;
     c(11) <= g(11) or (a(11) and g(10)) or (a(11) and a(10) and g(9)) or (a(11) and a(10) and a(9)  and g(8)) or (a(11) and a(10) and a(9) and a(8) and g(7)) or (a(11) and a(10) and a(9) and a(8) and a(7)    
                 and g(6)) or (a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and g(5)) or (a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and a(5) and g(4)) or (a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and g(3)) or (a(11) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3)   and g(2)) or (a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y10 or x11;
     c(12) <= g(12) or (a(12) and g(11)) or (a(12) and a(11) and g(10)) or (a(12) and a(11) and a(10)   and g(9)) or (a(12) and a(11) and a(10) and a(9) and g(8)) or (a(11) and a(10) and a(9) and a(8)    
                 and g(7)) or (a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and g(6)) or (a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and g(5)) or (a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and g(4)) or (a(12) and a(11) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4)  and g(3)) or (a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and g(2)) or (a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y11 or x12;
     c(13) <= g(13) or (a(13) and g(12)) or (a(13) and a(12) and g(11)) or (a(13) and a(12) and a(11) and g(10)) or (a(13) and a(12) and a(11) and a(10) and g(9)) or (a(13) and a(11) and a(10) and a(9)    
                 and g(8)) or (a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and g(7)) or (a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and g(6)) or (a(13) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                  g(5)) or (a(13) and a(12) and a(11) and a(9) and a(8) and a(7) and a(6) and
                 a(5)  and g(4)) or (a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and g(3)) or (a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and g(2)) or(a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y12 or x13;
     c(14) <= g(14) or (a(14) and g(13)) or (a(14) and a(13) and g(12)) or (a(14) and a(13) and a(12) and g(11)) or (a(14) and a(13) and a(12) and a(11) and g(10)) or (a(14) and a(13) and a(11) and a(10)     
                 and g(9)) or (a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and g(8)) or (a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and g(7)) or (a(14) and a(13) and a(11) and a(10) and a(9) and a(8) and a(7) and 
                  g(6)) or (a(14) and a(13) and a(12) and a(11) and a(9) and a(8) and a(7) and a(6) and
                  g(5)) or (a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and g(4)) or (a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and g(3)) or(a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and g(2)) or (a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y13 or x14;
     c(15) <= g(15) or (a(15) and g(14)) or (a(15) and a(14) and g(13)) or (a(15) and a(14) and a(13) and g(12)) or (a(15) and a(14) and a(13) and a(12) and g(11)) or (a(15) and a(14) and a(13) and a(11)     
                 and g(10)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and g(9)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and g(8)) or (a(15) and a(14) and a(13) and a(11) and a(10) and a(9) and a(8) and
                  g(7)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(9) and a(8) and a(7) and
                  g(6)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                  g(5)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and g(4)) or(a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and g(3)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and g(2)) or (a(15) and a(14) and a(13) and a(12) and a(11) and a(10) and a(9) and a(8) and a(7) and a(6) and
                 a(5) and a(4) and a(3) and a(2) and g(1)) or y14 or x15;                   

END behavioral;	
------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

ENTITY cla_16_32 IS
PORT ( din1, din2 : in STD_LOGIC_VECTOR(31 downto 0);
       dout : out STD_LOGIC_VECTOR(31 downto 0));
END cla_16_32;	  

ARCHITECTURE behavioral OF cla_16_32 IS
signal c: std_logic_vector(1 downto 0);


component cla_16 IS
PORT ( din1, din2 : in STD_LOGIC_VECTOR(15 downto 0);
      c0 : in STD_LOGIC;
      c16 : out STD_LOGIC;
	    dout : out STD_LOGIC_VECTOR(15 downto 0));
END component;

BEGIN
	

cla_16_1 : cla_16 
      PORT map( din1(15 downto 0), din2(15 downto 0), '0' , c(0) ,  dout(15 downto 0) );

cla_16_2 : cla_16 
      PORT map( din1(31 downto 16), din2(31 downto 16), c(0) , c(1) ,  dout(31 downto 16) );


END behavioral;	 
------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY cla_16 IS
PORT ( din1, din2 : in STD_LOGIC_VECTOR(15 downto 0);
      c0 : in STD_LOGIC;
      c16 : out STD_LOGIC;
	    dout : out STD_LOGIC_VECTOR(15 downto 0));
END cla_16;	  

ARCHITECTURE behavioral OF cla_16 IS
signal c, P, G, A : std_logic_vector(15 downto 0);

component GAP_16 IS
PORT ( din1, din2 : in STD_LOGIC_VECTOR(15 downto 0);
       P,G, A : out STD_LOGIC_VECTOR(15 downto 0));
END component;

component CLG_16 IS
PORT ( P,G, A : in STD_LOGIC_VECTOR(15 downto 0);
      c0 : in std_logic;
       C : out STD_LOGIC_VECTOR(15 downto 0));
END component;


BEGIN
	
 mu_gap : GAP_16 
  PORT MAP( din1, din2, 
       P, G, A );
       
MY_CLG : CLG_16 
  PORT MAP( P,G, A,
      c0 ,
       C );


c16 <= C(15);
dout(0) <= p(0) xor c0;
dout(15 downto 1) <= p(15 downto 1) xor c(14 downto 0);


END behavioral;	
------------------------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY GAP_16 IS
PORT ( din1, din2 : in STD_LOGIC_VECTOR(15 downto 0);
       P,G, A : out STD_LOGIC_VECTOR(15 downto 0));
END GAP_16;	  

ARCHITECTURE behavioral OF GAP_16 IS
BEGIN
	
p <= din1 xor din2;
G <=  din1 and din2;
a <= din1 or din2;

END behavioral;
------------------------------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity single_port_RAM is
  generic ( n : integer := 15;
			addr_width : integer := 4 ;
			row : integer := 4 
			);
  port(
    clk: in std_logic;
    we : in std_logic;
    addr : in std_logic_vector(addr_width downto 0);
    din : in std_logic_vector(n downto 0);
    dout : out std_logic_vector(n downto 0)
    );
end single_port_RAM;

architecture arch of single_port_RAM is
 -- type ram_type is array (2**addr_width-1 downto 0) of std_logic_vector (15 downto 0);
 type ram_type is array (row downto 0) of std_logic_vector (n downto 0);
 signal ram_single_port : ram_type := (others => (others =>'0'));
begin
  process(clk)
  begin 
    if (clk'event and clk='1') then
      if (we='1') then 
        ram_single_port(to_integer(unsigned(addr))) <= din;
	  else 
  		dout<=ram_single_port(to_integer(unsigned(addr)));
      end if;
  end if;
  end process;


end arch;
--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
    generic(
        addr_col  : integer := 10; -- required bits to store 16 elements
		col : integer := 1023;
        addr_row  : integer := 4; -- required bits to store 16 elements
		row : integer :=12
        );
	port(
		addr_c : in std_logic_vector(addr_col downto 0);
		addr_r : in std_logic_vector(addr_row downto 0);
		data : out std_logic_vector(19 downto 0)
	);
end ROM;
	
architecture arch of ROM is

    type rom_type is array (col downto 0) of std_logic_vector(19 downto 0);
	type map1_rom is array (row downto 0) of rom_type;
    signal weight_ROM : map1_rom ; --:= ( others =>(others => (others =>'0')));

	begin
		weight_ROM(0) <= (
		 "01001010101101011010", "11001110101100111000", "01000001100100101100", "11010010001101010111", "01001110001011101010", "11000110110100110111", "11010110000100000101", "00110110011100101000", "01000110000011100111", "11000010011100011010", "10101010001100011100", "11011110011100000111", "10111010010100000100", "01001010011100100111", "10111110000011111000", "11011010100100010110", "11001111000011100111", "11000010010100011001", "11000010010100000111", "01001111010100010101", "01011101110101011000", "00110001110100100111", "11000110011100110111", "00110110010101000101", "01100101110100110100", "11000001111101010101", "01000010001100111000", "01010001110101011001", "10111010111011110101", "10111010010011101001", "11000010010100100111", "11010010000011000100", "01000010000111110101", "11011110011101100101", "01001110011101011000", "01000111100100101000", "00110010011101010110", "11000110011111000100", "10110110011100100100", "10111001111100100101", "00111001111100011001", "11010110101100110111", "10111101100011101111", "11000101111100011000", "01010010111100101011", "01010010100110000110", "01001010000011100101", "01001110010100001100", "00101011000011111000", "11001010000011101010",
		 "11101110000100011000", "11000110101100101000", "11001001111100011000", "00111010001011100101", "01001110010100110100", "01111110010100000110", "10111110000011110110", "10111110011100001001", "11001110001100110110", "10110010010100101000", "00110110011100010100", "01000010000101111001", "01001001110110110100", "01001010010100000111", "00111010000100010110", "01010110110101110111", "10011110011110010111", "11010001111100110011", "10111101101011111011", "11000010011101011000", "01011110000101001000", "00111010110100000100", "01000110001100000111", "10111010101101011001", "01111111100100110110", "11110010001100101010", "01001010100111111000", "01000010001101111011", "11010010011101010111", "11011110011100011000", "01000001110101011011", "11011010011011101100", "00101010111011111011", "11000110000100101010", "10111110010110000111", "01100010000011111000", "11000010101100100011", "01011010110100001000", "01001101111101110111", "01010110001011111000", "10111010001100111000", "01001110111100100110", "01001101110100000111", "01000110010100110111", "11000001110100010111", "10110010000100000111", "10110010100101101000", "10111001110100100110", "01000010010110000111", "00111101111101000100",
		 "11001010011101110100", "01010110010111011000", "11000010110011111000", "01000110010100010100", "00111010001100001010", "01010101110100010111", "01000110000101011000", "11001110110100000111", "01000010000100010110", "01010110001100000100", "01010110100101101000", "11011101111101010111", "01001010101110001000", "10111110011100001100", "11000101111011111100", "00111111001100010111", "11001110110101111001", "01001010000100001001", "10110010001100100111", "01001110011100001011", "11010110011100001000", "01000010111100010110", "11000110010100001010", "01010010001011111010", "01010101110100010110", "01000110100100000101", "10110101110100001000", "10110110110110101000", "10111010000100000110", "00101010000110000111", "10111110011011110100", "11000010100100010100", "01001110010101100111", "00111010100100101001", "00100101100011001001", "10110101100100100111", "11000110010100111000", "10110110000101010111", "11000001111100010111", "00111110000101111010", "11000010010100110101", "00111010001100000110", "11000010000101111100", "11000010010110000110", "11011010011101111000", "11000110001101000111", "00110010011011000011", "11000101110101010101", "10111111100011110111", "00111110010100101000",
		 "01000110001011101011", "10111001110011101000", "10111101110101110111", "00111110010100010110", "01011101110100100110", "01011110011011110111", "00111110000111111000", "00111110010100001001", "01000010010100011001", "11000110001101100110", "01100010101100011000", "01000010000100101010", "00111110001100100111", "01010110010100101010", "01001110011101010100", "10110011100101110111", "01000001111011111001", "10101101111100011001", "10111001111011110110", "10111110001101010110", "00111010011101010111", "00110110001100001000", "01000110011100011001", "11010110011011111001", "01010010000100101000", "10100101110110001010", "00110011000011111000", "01001010000100110100", "00110001110011000110", "10111010100011101001", "11000001111100110101", "01001110001110111001", "10111010000100000111", "01000011110100110101", "11001110000100010110", "11000001110101011000", "11100101110101101101", "01010010000101100101", "10111101100100011000", "11000110101011110111", "01001101110011010101", "01001010010100100100", "01001110001011111000", "01010110000100100111", "01000110010110010100", "10111110011100000110", "11010011110010100011", "11000110011100101010", "01000001111110001000", "01011110110101010101",
		 "11001110011101101100", "01010010111011100110", "01001110010101010111", "11010010001100000111", "10110010111100110101", "11001110101100100110", "01001010011100101011", "10101110000100110111", "10110001110100101010", "01001110111101101001", "00101001111100001011", "11000110011011100111", "11000010010101010101", "01110110101011111010", "10100010010111001010", "01001110100100110110", "11000010000101111000", "01101110001100110110", "11011110110101110101", "10111010001101001001", "01011010011100111000", "01001110101100100101", "11001110111111010011", "10110001110100001001", "10111010001100010101", "10101110001100010101", "10101010010100101001", "00110001101101001000", "11000110100101101000", "11001010010100101010", "10110010011110101000", "01000010011100001110", "11000110010100010111", "11001110011100011000", "01001110010011110111", "11001110100101110111", "11000010011100101001", "00110010011110001001", "01011111100101001011", "00111011011100000110", "00111110111100000101", "11000110011100010110", "10110010001100010110", "01010010010100110111", "11000111010100101001", "00111010101100100110", "11010110000101110110", "10111110000011111000", "00111010000110100110", "01000110011100001000",
		 "00111001111100001010", "10110101111100111010", "01000011001100001000", "10110110010110100111", "00110001100100101001", "11001110000110010111", "01111010000100111000", "11001010110100111001", "00101101100100101010", "00111110000010110111", "10111010101100111001", "11000101111011110111", "00110111011101101010", "10111010010011111110", "10111010111100111010", "11010110110011101010", "01011010101101010101", "11001110100101000101", "01010010010100011000", "01000010010100110110", "01000010001100010110", "01101110010011100101", "00110010010101001000", "11001010000100010101", "11001110010101101001", "11001110001111010111", "00110010001100101001", "00101010101101001000", "11000110000011110101", "01001110001101000100", "10111110001100101010", "01000010000100010110", "01001110001100010101", "01100010010100101001", "01000010010100001001", "01000010010100001011", "10111110011101001101", "00111001110100010110", "00111010011100010111", "10111110011100100110", "01010010001100101010", "10111010101100111010", "11001111000100001001", "11101010011100101100", "11001110001101000110", "01101101111011100011", "01001101110101011100", "00110110101011101000", "11101010001100001100", "00101110001101000101",
		 "01001110000100010110", "01001010001011110110", "10101110001101010110", "01001001110100100110", "01000110001101110110", "10101110001100011000", "00111010000011101001", "00111110111100101001", "11000101110101101000", "00111001110110001000", "10101010000100000111", "11000010010100101000", "01101010111100111010", "10101010100101000110", "10111010010100101001", "10110001111101000101", "00111111000110000110", "10110110101100000111", "00111101110101101000", "10111001110110011000", "11000101100101001011", "01000010101100000101", "00110011001110010110", "10110010010101110111", "01000110001100010111", "01001110010100010101", "11000010000100111001", "10111010000100000110", "00110101101100110100", "01010010111100010111", "10100110001100111001", "01000110000100111001", "00110110000100000111", "10111110111100001010", "01010111010100010110", "01000011000100010111", "10111010000100010101", "11100010001100011000", "01001110000100100111", "11000110011011010110", "01001110110100000100", "00110110011011110101", "11000110011100101001", "01000010100101000111", "11001110010100000101", "11001110001100011000", "10101001110100000110", "10111010100100101000", "11001001111100010110", "00111101110100010101", 
		 "11001010110100110111", "10100001001111000111", "00110101011110001001", "11000001111101010110", "01000110111100000110", "10101101110101001000", "01000010000100000111", "10110110000100011110", "00110010011100100110", "10100010000100001010", "10100010101101101001", "01111110011100011000", "10100001111101100100", "01000001111011100111", "01001010010100000111", "01001110010101010110", "10110110001100100110", "00100110100011010110", "10111110000100000110", "01000110010100010011", "11011110010100110111", "10110010001101001001", "11001110111100011000", "10111110011100010101", "01000010001101010101", "10111110000101100111", "01001110000100011010", "00111010001100111000", "10110110110100110011", "00111001111100111001", "11001010010011111010", "00111110110100000100", "00111010101101100010", "10111010000101010011", "10110001110100110110", "01000101101101010101", "10101101000101000111", "01001001111100000111", "00111001111100100111", "01000010100101100100", "00101001101100001100", "11001010011101010100", "10100101001100101000", "00111010000100010111", "11000110010110000111", "01000010000100101000", "11000101110111111000", "01010001111110001001", "00011010000100100110", "10110010000100001000",
		 "01000011100011110111", "10111001111100111000", "01010010011100001100", "00110001111100110110", "00111101110101001000", "00101010100011000110", "01001010000011110100", "10110001110100010111", "11000010011100110110", "10110010010100000111", "00110010100100110011", "00111101110100110110", "11011101110100001001", "10110110011100011000", "11001001110100010110", "01010010101101010110", "10101101110011100111", "00111101111110100111", "00011001111100011101", "10110110010100110101", "00101001111100011001", "10110001101011100101", "10101110001100000110", "00101110000100000111", "00110010001101010110", "01010101111100010110", "00111110010100110100", "01100010011100101001", "10110111001101000110", "01010011001011000110", "01001110001100001100", "10110110100011111010", "00100101111100001010", "01000110010100101000", "10111010010011110101", "00111010001011001000", "00111110101101000101", "01010111000101011000", "10110010110100100101", "10110010000011001000", "10110010011011110111", "00110010010100000100", "11000101100101001010", "11011110001101110100", "00111110010101001000", "00110001110100100110", "10110010000101010110", "10111110101011010110", "11101110100100111100", "00101001110100000100",
		 "00101110000100100101", "00101110110101111010", "10101001110011000101", "00111010111100110100", "00110001110100011000", "10111101100100110100", "01100010000100110100", "00110010100101000100", "01010110001100110110", "01000001110011000101", "01001001111100000101", "11001010100100100111", "11001010011101010110", "10110101111011000111", "11000110011100010111", "01001010100100011000", "00111110011011000101", "10101010010101001001", "10110110010011010111", "10110101011100001000", "10101110000101010111", "00110110101100100011", "00110101111100000101", "01001010010100111001", "00111010001100000011", "10101010001011100100", "00110010000100100110", "11001101011101110110", "10101101111011110110", "10110101101100001001", "11010010101011110100", "11001110000100110011", "01000110011101011000", "10100101110011100110", "10111001000011100101", "01010101100011101001", "10101101110100001000", "10101010100100100101", "10100001011101010101", "01100110001100100100", "10111001101100000111", "10111001011011100101", "00011001100100010101", "00111110101011100111", "01111010001100010110", "11001010100110100101", "00110101110010100111", "11001010011101010110", "10101010000011001000", "10110110001100100110",
		 "01001010011011111001", "01001001011100100110", "10111001110100010111", "00111010011101100111", "00110010000011100011", "00110101101100110111", "11011110110011110101", "01001001100100000100", "00111111000100101000", "10100110000100011000", "11000001111011010101", "01000010000100100011", "11001010101011100111", "01001110101011111001", "00111001111011010101", "10111011100100011010", "11000101110011101001", "00111101100010101001", "10110010000101011000", "01010001100100000101", "10111010010011101000", "00101010000100010111", "10110110101100110101", "11000110001010101101", "10111111000100100110", "10011101111101001001", "10110101110011101000", "10110110100100010110", "10100110001011100111", "00110010000100000110", "00111001110101010011", "01001101110100000111", "10100010101100111010", "11011010001011000011", "10100011010100101010", "10110010001011001010", "01010010000011111001", "10110010000011000111", "10100101010101110110", "00110010001100010110", "11000001110011010100", "11100111100100100110", "00101110011100100111", "11000001111011010011", "10110001100010010110", "10101010001011100101", "10101001110011101001", "10110010001100100111", "01000010000101100110", "00110010011011010100",
		 "10111110001100111001", "01000010100011100110", "10101001111011000110", "00111110001100010011", "10111110010101010110", "00110010001011100011", "10111010001101101000", "10110010000011101001", "10100010101010101001", "10111001110101111001", "10110001010011111000", "10100110010011000110", "11011010001100101010", "00111110001100001000", "11000010100101001000", "01001110001100010101", "00101110011100110111", "11011001111100110101", "11000111000101010101", "01100010000011111001", "01000010010100000110", "01001010010100000110", "11001010111100110111", "10110001110011011000", "10111001011100010101", "10110110001100100101", "10101101010100011001", "00100110100100000110", "11000101111110001000", "11001010101011110111", "10110010011011101000", "01111010001100111010", "10110110011011110111", "11010101110110110111", "01010101100100010111", "10111110011011010110", "00101010010011101001", "00100110001101011011", "10110101100100110111", "01111010110100100110", "00111010000100000111", "01001010001100110101", "10111010111011110101", "11011110001100010101", "11001010100101001010", "11000110111100110101", "10110010100100100111", "10101010010100011001", "01101001111011100111", "10111010111101010111",
		 "10111101100101011100", "10100001010101111010", "10110101111100010111", "00100010001100111001", "00100001010011100111", "00110010011110000101", "11001110010100011001", "11000110010100101000", "00010101110100000101", "10101101100010101001", "11000111010101100111", "10110001110011001000", "10101110011100001010", "10100010100011000110", "10110101010100110110", "01000101011011011001", "00110001101011000110", "10111101101100010110", "10110110011100100111", "10110010001101010110", "00111010001100110110", "00110010101100100111", "11010010000011000110", "10110001010011101001", "10110110001011100101", "10111101111100101011", "00101010010011100111", "10110001101101000101", "00111010011100000101", "10100110101101010011", "11001010101100010110", "11000110100100110100", "10111110010101000100", "11000010001100101001", "00101110001011110101", "00111010000101001000", "01001110110100111001", "10110011000110010111", "00110001110101100100", "10101010010100100111", "10111101101101010110", "00101010011110011000", "11001010011101011000", "10110010000110000110", "10111010010101000110", "10101110101100100100", "10111010011110111011", "00111010100011100111", "00111110001100000111", "10111010001011100011",
		 "01100010101011110100", "01011010010110110111", "00110011111011010101", "00100110000011100110", "00110010001101110111", "10100101110101001000", "10111111001100000100", "00101010001011100110", "10111101100100000111", "10111101110100001001", "10011110010110100111", "10111111011011010111", "10111110010100010111", "00110010110100000101", "01010001110100011001", "00111001111011100101", "01001010010011110101", "00111110100100000011", "00101001100100100111", "10111010000100001000", "01010010010100011010", "00101110001100000101", "11000101110101110110", "00101001011100010100", "10111010011100000101", "01000010101100110100", "10110010011100010110", "01000010010011110111", "00110001010011001000", "01001110011100110111", "10101101111100000110", "01001010101100110101", "10101111010100010111", "10111001111101100111", "11001001110011110110", "00111010100011110011", "10101110010100110101", "01001110000100001000", "10111010000011110101", "10101110000010111000", "01001010000011100110", "11011110001100010110", "10101010010100001010", "00111010001011110111", "01000110100010110101", "00101001110010100110", "00101110101100100101", "10101110001110011010", "10111110010110110110", "00100010011011001000",
		 "11000110101100001000", "11000010001101000111", "00111001101011101001", "00111110011011100111", "01111010011011001000", "10111010001100101001", "00110110000100001001", "10110101101101011000", "01000010000100011001", "00011010100011000111", "10111110101101001000", "10111010001101000100", "00110001111011100101", "00111001111100101100", "01001110110110000101", "10111011011100000101", "00110110011011010101", "00110010011110010101", "00111010010100010110", "01011101110101011000", "01000010001011100110", "00100001011100010101", "11000101110100010110", "10111110001100000111", "01000001000011100100", "00111110000100110110", "00111110000100010110", "11001110101100000101", "10111010001100110100", "10101101111101000111", "01001010010100011000", "01011010000011110110", "01000010010100000100", "00111110011100010110", "11000001111100101000", "00110110100010111000", "10101101011101001001", "00110001111011100100", "11001010001011100011", "10110101110100110110", "01001110000101011000", "10111110000011100101", "11000101110100000111", "00111001111101011000", "11000110000110000111", "01010011110100000011", "01000110101100100101", "11100010111101110110", "01000010110100100111", "10111010000100011001",
		 "01011101111011110110", "10111101110100101010", "11100001111011111001", "10111110001101010101", "00111001110101000100", "00110110111100000100", "01111010000011110100", "11001010000100000011", "01000110000100010110", "01100110100011100111", "00111101111100000100", "11011010101100111001", "01001101100101000110", "11000010010100001000", "10111110011100110110", "01010010101101010110", "10011101010100111110", "10110110000100110011", "01000101111100101000", "00111110101100011000", "00111110100101010110", "10101010000011110110", "11001110000100111000", "10110101110101001001", "00101001110100110111", "01000101110101011000", "01010110000011011001", "01001110010011100111", "01000010000100000101", "01010110010100011000", "10111010100101100110", "11011110011100110111", "10101011011010101001", "11010110011100110111", "00110110111101000100", "00110110111010100111", "10111101110100000100", "01000011000101000101", "10111010011101010110", "00100010101100101000", "10110110011011001000", "10110001111100100010", "11001010010100101000", "01000110010100110111", "11001110101100110111", "10110001111010100100", "00101001110100010110", "01001110011011100101", "11001010000101001000", "00101010011100100101",
		 "00110010101101010110", "10111010010100000110", "00101010010111101000", "10101010001100000100", "11000010011100100111", "10111101110011111000", "11000001110100110101", "10110110000100010101", "01001010010100010111", "00111001100011000110", "00110001110101000101", "11000011101011110111", "01001110110100011000", "10111110001101101000", "00110011111110011000", "00110010000100100110", "11000111101100000101", "11010010000100001000", "00110110010011001010", "00100010001100001000", "10111110101100011001", "01000110101011010101", "10111010011011101111", "11000011000101011010", "10111010011100000100", "10110011101100100111", "00011101111100001000", "01000010000100000101", "00101010011100000101", "10110101111010101011", "01000010010011110101", "10111111000101010101", "00101010100100011000", "10100010010011110101", "10110001110010100101", "10111101110011101010", "01010101110011001000", "10110110010110010110", "10110001110111101000", "11000110001100010110", "11000101111011100101", "10101001011011000100", "00101001110011100011", "01000110000100010101", "11001010101100000111", "10111010001110010111", "11001001110011010110", "10111101110100010101", "11000110011100010101", "11001010000100110100",
		 "01010110010101100111", "10101101111100000111", "11000110111100101000", "01000010100100000101", "10111110100100100100", "11011110010101001000", "01000010011101001010", "10110110000011000101", "11001110101101001001", "10101010001100111001", "11010010011100010011", "01111101111101100100", "00101001101100000111", "10111101110100111001", "00111010000100010101", "10110101100110010111", "11000110100011110111", "00011101100010101000", "00100110011101010100", "10111001101110000011", "10101010000100110100", "10100110000011111000", "11001110011100010011", "11000010001011101000", "10111110000100110110", "11000010100100101010", "00101101111011011000", "10101110010100000110", "10110010000100010110", "00011001100011000110", "01000010010110000111", "11001101110101010110", "10101010011100101001", "00110001101011110011", "00110110010011110111", "01000110011101010111", "11010001101100111000", "10110110010100000110", "00101010001101100101", "01011110001100010100", "00110110000010100100", "00111011000100000100", "00100101011100001000", "01001010010101010100", "01000101110011110111", "10101110001100000100", "00110110011100000100", "10110011010011011001", "10111110010101100111", "01000101110100000101",
		 "00101010001100100101", "11001010000011110110", "11000010010100101001", "00111010000011110101", "10111010010100010110", "01010010000101010110", "01000010001100111001", "10111110110100111011", "00110111000011110111", "11000010010101011010", "00110001111100101001", "10101001110010110101", "01001011010111110100", "01001101111011101010", "00110110100011100111", "11001101110100110100", "00110110010100111100", "00111110010100001000", "11011010011101010110", "01010010101100101000", "11011010101100110110", "11010110001100011001", "01000110010011110101", "01000010001011101000", "10111010000100010101", "10101010101011110110", "00100110000100011010", "10110101011011000110", "10111101100110010110", "11001010011100001000", "01001001110101000110", "00111010000100000111", "10101110000100111010", "10110010000100111010", "10110101100011110101", "01000011111100110101", "11000001100100001000", "10110001111110001000", "10111110010100111000", "00110010000100000110", "00110001100100110110", "01010101111101010101", "00111001001011100100", "10111110011011010111", "01001110010100101001", "01000010001110000110", "10101101101101010100", "01001110011110000111", "11000110011011001001", "01001010000110011000",
		 "10111101111100011011", "00101110000110001000", "01011001111011101010", "00101010000110100101", "00100011100011101000", "11000011000100010111", "00111110001011001000", "11000110101101101001", "00101101011100110101", "00100101001011011001", "00111010001100101000", "10111001110011101010", "10101001110101001000", "10111010000011101000", "10101110000100010101", "00110101110111001000", "01011001101011100100", "00110010001100100110", "10101110010100100111", "10111110001101110101", "10110110111100100101", "10111110101100010100", "10110101101101000110", "10111001111100000100", "00110110001011000101", "11000010000011101001", "10110110010100111000", "10110101100100111010", "11001110011100000100", "01111110010111110111", "11011010000101000111", "00111001111100010110", "01001010000100010111", "11001010001100111001", "10101110100111100111", "01000110010100000101", "11010110000100111000", "00111010000100101111", "11000001110100110101", "10111001111100100101", "01111110001100111001", "10101110000101100111", "01000110111011100111", "11011110000100000110", "11000010011100100101", "10101101111100100101", "01011010000100101010", "10101110011101000110", "01001010111100010111", "00111001111100000011",
		 "10110110101100101010", "10101101111101000111", "01000110000011101000", "00111001111011100111", "01010110001100011001", "10100101111100100101", "00110001110100010100", "11000101110101011011", "00101010000100101001", "11010101101100101001", "11000001100111100111", "11000110011100110111", "01001001111100110111", "01000001110100111010", "00111110101011110110", "10111110001100011010", "11010010011100110100", "01000001110100010110", "01000001110100011000", "11010111011100110110", "00110010111010101001", "10111101110100111010", "01000010000011001000", "00111001111011100111");
		weight_ROM(1) <= (
		 "01000110011110001001", "01001010101101001001", "11001010010100011010", "11000010000100001001", "11010010001100101001", "01001011011100111000", "01001010011100111011", "01001010001101111000", "10111010011100111001", "00111110101110101001", "10111010010101011011", "11001010011100011001", "11000010000100001101", "01100011100100011000", "11001110000100011000", "11000010000100101010", "11000110110110000111", "11000010010100101001", "11001010010100001011", "01001010001100101001", "01001010011101001111", "11000010011100001100", "01001010100101011110", "01111110001100001100", "01001110010101101001", "11101110000101110111", "10111110010100111000", "01001010100101101001", "01010010010100001000", "11000110101100111101", "01000010010101101001", "01010110101100101100", "01000110010100101010", "00111110110100101010", "11101010011101001000", "11000110000100111001", "00111010010100101010", "11000110110100001001", "01010010100101001000", "11000110010100001001", "01000111000101101000", "01001110100100111001", "11001110000100101010", "11011110001100011000", "11010010000101001000", "11000010011100101000", "01000110010100111000", "11001110000111110111", "01000010011100101101", "11000010111100001000",
		 "11010110010100011001", "01000110001100001011", "01001110000100111000", "01100010010100001001", "11000010010100100111", "11010110100100010111", "10111101110100001011", "11010111010100101001", "11000110100101001010", "01000010010100101001", "11001010100110010111", "11010010011100011000", "00111010010100011011", "01001010011100101010", "01001110110100111000", "01001110010100111000", "01001001111101011010", "01001110100100111001", "01000110011100101000", "01000110001100100111", "01000010001100111001", "11010010001100101011", "01010010001100011011", "11010011000101011000", "11001101110011101110", "11010110100100011001", "11000010101100111001", "01010010010100001000", "01001010001101011000", "11010010111100001010", "01000010101100011001", "11010110010100011000", "10111011001100111101", "01000110011100101001", "01000010100100111011", "11000110000100111000", "11010010111100011001", "11000010011011101001", "11010110001100011010", "11000110000101101001", "01001010100111001010", "11000010110100001010", "11010110111100001000", "01000110001101011000", "01101010011011101001", "01011110100011111001", "11010110100101011001", "01000110000100101000", "11000110001100011001", "10111110001100101011",
		 "01000010000100111000", "11010110001100111000", "10111010000101001101", "01001010011110110110", "01011110010100111011", "11010110011101011010", "01001010001101101000", "11001110001100111000", "11000010101100101010", "11000111100100000111", "11000011000100101011", "11001110100100001011", "11010010100100001000", "01001110110101111001", "01000110001100000111", "01000110001101001000", "11010110001100001011", "10111010010101001001", "01000110011100011001", "01001010000100001001", "01000110000100111001", "11011010010100101001", "01010010100100011001", "01000110011100101001", "01010110000100011001", "11001110000100111001", "11000010000110111010", "01001110000100111000", "01001110011110111000", "11100110111100101000", "11001010001101011000", "11000110011100100111", "11000010000100101001", "11010110010100110111", "01111110010100011100", "01010110001011111000", "11010001110100011001", "01011110111100001001", "11001010011100000111", "01000110010100111000", "01010110001101011000", "11000110100100011001", "01000010000100001000", "11001011101110001010", "01000010000100111000", "01001110001100000111", "11000110100011111000", "01000110000100001100", "10111011111101011000", "01011010011100001001",
		 "11001010000111111001", "11001110010100101001", "11001110110100011011", "11011010010100111011", "01011110010100011000", "11010110101101011011", "01011110000100111001", "11001010100101001100", "10111010011101101010", "11000010011101111010", "00111001111101001000", "01001110111100011000", "11000110001101001001", "11001110011100111000", "01001010010100101000", "01001010001101001000", "01001110010100101000", "01001110000110001000", "01000010100101011011", "11001101111011100111", "01001110000100011100", "11000010000100001001", "11001110011100110111", "01000110010100011100", "00111010101101001110", "01010110000111101001", "01000010010100101100", "01010110001100001010", "10111011010101001001", "11100010001101010111", "11001010001100001001", "11001110100100110111", "01110010010101101001", "11000010001100001001", "11000110001100011000", "11000011000110001100", "11000010000101101001", "10111010101100101001", "11101010000100011001", "11010010110101011000", "00111010011100111001", "01010110000011100111", "11001110000110011010", "01000010010100011110", "11010011100101100111", "00111110101100011010", "01000010001101111000", "11000011111101101000", "11101111001110101010", "11001010000101011001",
		 "01000010010100011000", "11001111001100011011", "11001001110100001000", "01001110100100101000", "11000010001100000111", "11011110010100111001", "11100010000100011000", "00111011110100011101", "11010101111100011010", "11001110011100111001", "01001010001100101001", "01010010101110101011", "01000110101100101011", "10111010101011101010", "11010010000100101010", "01010110111100101000", "01010110001101111010", "11000010001100101010", "11001010010100011000", "11011011000100111100", "11010110001101001000", "11000010000100001010", "11001110100100011000", "01100010011101001001", "01010010010100101010", "01000010101100101001", "01000110010100011000", "01000110110100111001", "01000010001101001111", "01110010101100101000", "01001110011100101001", "01001010100101101001", "10111010010100101001", "11000010011100011000", "01001110000101011000", "11010001111100001011", "01100110001100001000", "11001110111100011001", "11010110010100011000", "00111010011110101001", "01010110010101001000", "11010010001100101111", "01000010101101101010", "01001110101100101000", "01011101110100111001", "01010110010101011000", "01000010000110011000", "01001101110100111001", "01000110011100011001", "11001001111100000111",
		 "11010010000100001001", "11000010001100101000", "01100010011101001100", "11000110000101001000", "01010111000101111001", "11000111011100111001", "11000110001011101001", "11010010010101011001", "11101110010110111001", "01001011111100011000", "11000010101100001010", "01011010000101101011", "01000110001100111010", "11001001111100101001", "11010010111011100111", "01001010011100111011", "11010010100101101001", "01000110001100111001", "01100010100100101001", "00111010010011101000", "01000110001100011001", "11101110011100001010", "11101010001110011001", "01010010101110110111", "01000010101110001010", "11001110000100101001", "11000110100101011010", "01000110111100111010", "01001010010101010111", "01010001110101001000", "10111110001100101010", "01000110011100011010", "11001010010100111010", "01001110100100011100", "00111110101100011001", "01001010000011101010", "11001110011100111001", "01001111011100001010", "11001010000110101000", "11001011000101001010", "01000110001100101000", "01011001111100011000", "10111110111101000111", "01111011001100001001", "01000110011100001000", "11001110011011101000", "01000110111100111100", "01111010011100111000", "01100010100011101001", "00111110001110001010",
		 "11001110010100101001", "00111110010100001010", "01011010100101011000", "11001101110101111001", "11000110101110001011", "01000110011100111001", "01010010011100001011", "01010010010100011010", "01100011000100010111", "01000001111100011010", "11101110110100001100", "01001010000100001100", "11100010011100101010", "01101110001101011001", "11000010010100101001", "11001110100100001001", "11000111000101011101", "11000011100100010111", "01010010000100101001", "01001010100100101001", "11000010001110110111", "01111010111110101001", "01100010011110001011", "01000010011100011001", "11000010011100011001", "11011110001100011000", "11000001110101101001", "11001010101100101001", "00111110110011111011", "00111110111100111011", "10111110000100001010", "11001010001100101000", "01101110000100110111", "01011110010100111010", "11010110100100001010", "01010010010100101010", "11000010010100001001", "01100010001100011000", "11011101111100001000", "11001010000100111101", "01011111001100001000", "01010110001110011000", "01000110000101101000", "11011110010101101000", "11011111000100001010", "00111010001100001011", "01001110010100001001", "01000110001100001001", "01111110101101101001", "00111101110100010101",
		 "01110101111100010111", "01001110100100101000", "00110101111111001000", "01001010000111011100", "01001110001100111000", "01011010010101011010", "11001110011100110101", "10110110000100111000", "00111110101100100111", "10110110011100111001", "10110001110100001010", "01110111000101101000", "11010001110110000111", "00111011000101011010", "01000110101101101000", "11100110001011101000", "11001110000100011010", "01011001111100111000", "11000110100110001001", "11000110010100010100", "10111101110111011001", "10111101111100101000", "01100110001100011001", "00111110000100101000", "11000101110100110110", "10111110000100111000", "11010110000100010111", "01000010000100111010", "11001010001101010110", "10111010001011101100", "01110110011100111000", "01011010000110100110", "11011110010101100100", "01000110010100110101", "01000010001011101001", "00110110111100110110", "10100101100101000110", "01000010001011110111", "00110111000111000100", "11010010011100001000", "11000110100100011001", "01001011000110011000", "01000101111100001001", "11010010000100011000", "01001110000101011010", "11001110010011111110", "00111010011100010101", "11000011010100011001", "00100110010110111010", "11010110011100101000",
		 "01001010001101111001", "10111010100011111010", "11000010000100100110", "10111110101100111000", "11000010001100011001", "00111110001101000101", "11010110000100010111", "01000010010101100100", "01000110101101010111", "11000111101101001001", "01000110011101010100", "01010010100100111000", "10111110111110000110", "01000010010101111001", "10110110001100101001", "11010110011110101011", "11000101100101011001", "11010110000100110111", "00101010001101000111", "01000010000101101011", "01000110111100001010", "11000111011011100110", "11100101111100001000", "00111010000100101001", "01000010011100010110", "01001010000100011110", "11000010100111011000", "11010011001101011001", "11011010010100011010", "01001010111100010110", "01100110001100101000", "11001110010101001000", "00110101110100111001", "11000110001100101001", "11000111011100110110", "01011010001011111010", "00111110100110100110", "00110010101100111001", "01100010111100000110", "11000010111110010111", "10111010001011111001", "11001110001100100110", "11000010000101101000", "01001110001100110111", "01001110101100001001", "10111110010011101000", "00110010001101110110", "11000010101010110100", "11000010011100001010", "01000001111101100100",
		 "00101010100110000111", "11010110011101101000", "10110010010100001000", "11001110011100010100", "00111110011101101000", "01001010101100101001", "10111110101101110111", "01000010010100000111", "01000110001101011000", "01000110010110100110", "00111110010100001000", "11010010000101001010", "11000110001101001010", "11000010010100111000", "01000101110011101000", "01001110001011101000", "11011001111100000101", "11010010001101111100", "10111010010100011000", "00100110111101001000", "10111010110011110111", "01001110010101100101", "00111110010101111010", "01010110001011111000", "01000010011100100101", "10110110001100001000", "00101010000111011110", "11000101101101011001", "11011010001100010110", "01000110000100010111", "00111011001101011001", "11001010011101010100", "00111110000101011001", "10110010001100001001", "11000001001101000101", "01001110100101111000", "10101010110100101001", "01000010101101011000", "01001110001100001001", "01000010000100010110", "01001110001100010110", "10111001101101001000", "00100110100100110110", "00111110011100110101", "11010110110101011001", "11000111001110001000", "01000001110101010110", "01010110001101100110", "11000001110100000110", "01011010001100010101",
		 "11001010101011101111", "01001011011101001000", "10110101110110011000", "11000010100100010111", "01110111010100000101", "00111110011100101000", "01001110010111111010", "00111010011100101101", "10111010010100011010", "10111010010011101000", "01100110111101011001", "01011010101100100101", "10111110001100101000", "01010111101011101111", "11001010000101011000", "11000010000101101001", "01000110110110011010", "10111101100010101010", "01000110010100010101", "11011001111101000111", "01001110000101001000", "11000110001110001000", "11000110010100010110", "01000010010101011001", "10111110011101001111", "00101101110100011001", "01100111000100011001", "10110010010100100110", "11000110011100001110", "00101010001100110110", "11100010000100010101", "01111010010100110111", "01011110010100100111", "00111110000100100101", "11010110000100110101", "11100110011100001010", "01010010001100111000", "10111010100100111100", "00111010001100000110", "01010010001101010101", "11000110100011010011", "01100110001100100110", "11000110010100011001", "11010110101100010100", "11000110111100110110", "00111001110100100110", "10111110000010100111", "01001110001100001000", "11001111011011100111", "00110010010101110110",
		 "01001010011100011000", "11011110100100100110", "11011110111011101001", "11001110011101101001", "11100110101011111001", "00110110000101000110", "01000010001100001001", "11001010111100100111", "10101110100011111000", "01001110011101001000", "00110010100011100111", "11010110011100001000", "01001101110101010110", "10111011001100111000", "11010110010100001000", "01011110010100011001", "10110110000100111000", "01011101110100100111", "11000110101101010101", "01001101110100011000", "11000110101011101001", "01001010001101111000", "01010110011100100110", "00110101111100011000", "10111110000110100111", "11000010011100100111", "11001101110100110111", "00100010010100100111", "01000011001100000111", "11000010011100110111", "10110110001100010111", "11001001110011101001", "01001110000101101101", "10111001110100001000", "10101101111110010111", "11000010000100110110", "11011110000100000111", "10111010010100001001", "10111110101011111000", "11010110011110110101", "00111010000101001000", "11101011001100111000", "00110010000100101000", "11001110011101001000", "01001110010100111001", "10111010000100110110", "10111110001100101000", "10111001110111011010", "01010010010110011000", "01000001110100011011",
		 "11011010011100011100", "10111101111100101001", "01011010100101000111", "00110011000100001001", "01000010000101011010", "01010010101100110110", "11011110000101001010", "01001010100100101010", "00011110011101100110", "00110010010010101000", "01101110100111000111", "10111011000011111000", "10110010101100011010", "01010110000100000111", "01001011001101011001", "11001101111101011010", "00111010010100000100", "01000010000100100111", "11000110011100100111", "11010110010100010101", "01000110110011100100", "01000010001100101101", "01000110010100010110", "11001010110011110110", "11000101111011100110", "01000110010100110111", "01000010000011100111", "10111110001100000111", "11001110101100000110", "10111110111011110100", "01111010011011100111", "11010010000100110100", "01011010101011110111", "11001110001100011011", "01000110010110011000", "11001110001011110111", "11010010011011111000", "01000111000100000111", "01000010011100100111", "10111010100100000101", "11001110100100111001", "11000110011110011000", "01110010000011111001", "11000010001100010111", "00111010101101001000", "10111110010100100101", "01001110001101101010", "10101110001110010110", "01010101111100010111", "11001110000101100110",
		 "11000110000100111011", "11000010010101110110", "01000010000101011000", "01000110010100011000", "01011010000100000111", "10101010100100001000", "01010010100011100111", "00110010001100100110", "01110010000101001001", "10111110001100111000", "10101110101100001011", "01000110110100001000", "11010010010101011000", "10111101110100001010", "01001001111100111001", "00101010011100111001", "11000101110011110101", "00101010100011000101", "00110001110101011010", "10110110011100101010", "11000110011101001100", "00101110010111100111", "01001010010101000110", "01000110011100000111", "10111010001100000111", "01011010010101110101", "10111001111100010110", "01000010001101011000", "01000010010100001000", "11010010101100010110", "10101101111101101000", "11000011110100100111", "11100010000100011001", "01000010101100101000", "01001110000100000110", "11000010100100010110", "11000010000100010110", "11011010011101111000", "10110101110101110011", "10110010010011110111", "11000010000101000100", "00110010010100110111", "00111110101100011000", "11001010101101101001", "11001110110100000110", "01001101110110111000", "00111110000100100111", "10110101111100010111", "00111110010100111100", "01001110111100100111", 
		 "01010110010100011010", "01000101111101101000", "10101101010101010111", "00110001111011111001", "00111011000100101000", "10101101100110100110", "01000011001100110110", "10111010010011111000", "00100001111101000101", "10110101110111000111", "01000110100011100111", "11000010001100010110", "11011011001100000110", "01010010000111000111", "01000010011100011001", "01010110110110011001", "01011010001011110101", "00110010100011101001", "01010010000100011000", "00111010010011111000", "11100001111011111001", "01010110011011101011", "01000110010011100110", "00101001101011000111", "00111110000011000110", "10110010011101000111", "11010010001100010100", "00101001110100110110", "01000010000100110101", "10110101110100011000", "11011110001100010110", "00110010000011100110", "10111110000100010110", "01000010000011110111", "10110110101100110111", "11000101110011011010", "00111110010100100111", "11011010011100001001", "00110010011011100110", "00110001110100000101", "00110010001100000111", "01000101111100101000", "00110110011100000110", "11000110100110100111", "11001001110100110111", "01001010010100000110", "00110001100110100110", "01000001110011111000", "01000001110100100111", "10111110001100001000",
		 "11000010010101011000", "10111110001100111000", "00110101111011111010", "00111010011100000111", "11010001111101010111", "00111110000011110100", "00101001110110101000", "10111101111011110101", "01000010011011000110", "10111010001011101000", "11000111000101010101", "01000110100011110111", "01000001100101111011", "10101110001100111000", "01011110100101101001", "11010011100101110111", "00101001000101000110", "01010010001100001011", "10111110100100001010", "11000010111100111000", "00111010010100110111", "01010010010011101001", "11010101110101010111", "10110101111110001011", "00110010010011110111", "11001010001011001001", "01001010001011010110", "01010110010100111001", "00111110010011111011", "11001110011100101001", "11000011110101000111", "10111101111100101000", "10110101111011100110", "11010110010011110111", "01000010001100011000", "11000110101101000110", "01100010010100000100", "01000111010100000110", "11001010011011111000", "11000010000011111001", "00110110000100111001", "11011010011110000101", "11000101111011100100", "01100010011100010101", "00110010001101010111", "00110010001011000101", "11000110011100001010", "01000001110100101000", "01000001111011110110", "10111010010100010101",
		 "01001010011101100111", "00111110110100110111", "11000001110011000110", "00110010110101001000", "10110010110011000111", "01100011011100101000", "11000010000101010111", "00101010000011110111", "00111010010100110101", "00101001110011100101", "11001010001101110101", "11001010000011110100", "00111110001100001000", "11001110000100100111", "10111101110101011001", "00111010101011111000", "01000010101100010110", "10110010000100000111", "11000110100100100111", "00111001111011001000", "10111011110100101101", "01000010001101010111", "01111110011100000111", "10101010001011101000", "00110001110011111100", "11001001111011111000", "00110110101011000110", "01000010001100110110", "01000001110011010111", "00111101101011100111", "11001010000100011001", "01000101110011001000", "00101010111100110111", "01000010010100010111", "11001110000100001000", "10111110010011101001", "10110001101101001010", "00111001101100000111", "10101110011011101001", "00111111001011100111", "01000101100011000101", "00110101111100010101", "00110001100100000111", "01000010011011100110", "01000010001011001001", "11001010110100011000", "00111010011011111000", "01010110101100100100", "01001110100011110100", "01001010000011100101",
		 "11001010011101011000", "00101110010011000110", "10111001100010100110", "10110111101011100110", "11000010000011010111", "10110101110100100110", "01000010111100111000", "10111010000100000111", "11010101111100001100", "11001110100011111001", "11010001101011100110", "01000010000100011000", "00110101101100000100", "10110101111011110111", "00111110001100010111", "10111110100100001000", "11000001110101001010", "11100010010011101011", "01010110101100000111", "11000110001101110111", "01010010001101110101", "10111010010100111000", "00110010101100010101", "11010110001011111001", "01000010000111011011", "10101010011011100110", "11000110011101001001", "11000010011100011001", "01001010000011100110", "10111110101100110110", "10111101110100010100", "11000110000011101001", "11000110100100111000", "01011101111011101111", "00110010000011100111", "10111001111011111000", "01000010011100000111", "01001010010100111000", "00101001100101100101", "11010110011100010110", "01001010000100011000", "01000010010100000101", "10111010001011101001", "10101010010100000111", "11000010001100011000", "01000010000011100111", "00111010100010100110", "11000011000100011010", "01000010000101000100", "00110011001011101000",
		 "11000110001100111000", "01000010000011100110", "11011101110100101111", "00110010000100000111", "00111101110100110111", "01010010000011110110", "00111010001100110111", "01001110010101011000", "10110101101100011011", "11000010010100001001", "11000010010101011010", "00111101111011101000", "10110110010100110100", "10111011001011110110", "10111001111100101001", "01010101110100010111", "00101010110011101001", "01001010100011100111", "01001110101100011001", "10111010001100110111", "11000010011100010110", "01010110111011101000", "11001010010011110101", "11001101010011111001", "00110110101011100111", "10110010000100100111", "11000101110011100110", "11001101111100010111", "01011010001011101000", "11001001111101010111", "01001101111100101010", "11000011010100001010", "10101110010100011000", "10110010100100101001", "00111010000011011011", "00111010000101100111", "10110110111100000111", "10101101110100001000", "11010101110011111011", "11011010010101110110", "00111010001011111011", "11000010000100010111", "00111111001011000110", "00110110000111100110", "10111010101101011000", "11000101111100111001", "00110110000011000111", "10110101110011101011", "00101001111011110100", "10111110001011001000",
		 "11000101110100111010", "10110110101011100111", "01001010001011001001", "10111001110101000110", "00101001110101100101", "11000010100101101111", "11011010010100001011", "10111010101100011001", "00110101111100100110", "10101101010011001000", "00111010000011111001", "01000110101111011000", "10111011000011101000", "10110110010100011000", "11010110001100111110", "11001010010100001001", "11000111001011011001", "10111101100011010100", "10110101110101111000", "01000110000011011000", "11010010010100010101", "10101110000100111001", "01000010010100011001", "01000101110011000111", "11000110101100110101", "10110011000011101000", "10110110011100001011", "00111101111011100111", "00111110101011100110", "01010101111011110110", "01001011011100100111", "11001110110100110110", "01000010111101011000", "11001010000011101000", "10110010011101000101", "01011001111011111000", "01000110100100111000", "10110011111011100101", "11000010001100110111", "11011010110011111000", "11000010011100101000", "10110101101100011000", "11001110110101011001", "01001010001100010101", "00110010100011100110", "11001110001011110110", "10110101111011010111", "01010011110011100101", "00111010010100100111", "00111001110011100110",
		 "11100101110101100101", "01000010011100010110", "11000010001100001101", "00111101110100100110", "11011001111011001001", "11010010001100000110", "00110101010100100111", "11100010010100111001", "10111101100101101000", "10111101111100011000", "10101110001101111001", "11000010000011000110", "10111110000110000110", "00111001111011100111", "10111010011100100101", "11001110101011110111", "11001010100011010111", "00111010000011110101", "11000010011101001000", "00110001111011100110", "00111010001100011000", "00101001111011111001", "10111101110100010110", "00111010001100010111"); 
		weight_ROM(2) <= (
		 "11000110011100011011", "00111110001011100110", "10110010011100001000", "00111010011100011000", "11001010011100011000", "10101010111011100110", "00111011100110010110", "10111011000011110111", "00100001110101000110", "10101101111110100111", "01011010000101100111", "01001101110100000111", "00111110011011100110", "01000001111100000111", "01000110001100010111", "11100010000011111011", "11001010011100011000", "11001010010101101111", "00110010011100011000", "11010010100100010110", "01001010001011101001", "10101110101100111000", "11010010011100101001", "00110001111011111000", "00111101110010101000", "10111110110100000111", "10111110010101010100", "00101001110100111000", "00111010000111111000", "10111010001100001000", "11001110011101110111", "01000001110011001000", "10110101100100011010", "11010001101101010110", "10111010100101110110", "11000001110100011001", "00110001110011100101", "11000001111100110110", "00110110101100000101", "00111010110011000110", "00110101101100001000", "00110101110011101000", "10110101101101000111", "01000110000100010110", "11011010001100010111", "01000001110100000111", "00101001110100111010", "00111001110011111000", "00110001110011001001", "11000110010100111100",
		 "00111010101100111000", "11001010100100101011", "01000010111011000101", "11010010001100000101", "01001001010011000111", "01001101110011001100", "00111001101100100110", "01000001101110000101", "01000110011011000111", "11000001101100000110", "11011001110110010111", "01000010000100010110", "11001001100011100101", "10101101101100101011", "00111010011100111000", "01001110000100010111", "00011001000011000110", "11000110000100110110", "10111110000100011001", "11001011011100100111", "10111110111110010110", "11011010101110011000", "11011110100100010101", "10101101110100101001", "00111001110100011000", "01011010101100101001", "10110110011100010100", "11001010000100011000", "01011110010100010111", "01011010011011100110", "01000110010101000101", "10111010010100011000", "01001101101011100110", "01010010001101100111", "01000010001101010110", "00111010001011000111", "00110001111101100101", "01000110000100111000", "11000110010100010101", "11001010100100011000", "00110001111011011000", "01101010110100000101", "11000011111011000101", "01000110011110001000", "01001001110101010111", "10101110111100001001", "11001010000100101000", "01000010011011010111", "00111010001100111000", "01010110110100010111",
		 "00110001110100100101", "00111110010011110111", "00110010010011001000", "01000010010011100110", "10100101110011010101", "10110010000011110110", "11000010001100010110", "00101110000011100110", "00111001110111110111", "00101010000011000110", "11001001110011011001", "11000110001100010101", "00111010011110001000", "01010101101100001001", "11000110000100001001", "01001111011100010110", "01000010011011001000", "10110001110100001000", "11000010010100000111", "01011101111100000111", "11000010000011101010", "00111111001011000111", "01001101100101011001", "10100110101011101001", "01000010000100100110", "01001110001100011100", "00101110111011000110", "00110010000011100110", "00111010100011010110", "00111010001101100111", "11001110100100010111", "00110110100011111000", "00101001110100111001", "10101110010101010111", "01001110100011101001", "11010001110100001000", "10101010011101001001", "00111001111100011000", "10110110100101001001", "00111010000101001001", "00111110010100100101", "01000001111011110110", "00100001110011101001", "11000010101100000101", "11000010011100001000", "01001010011110010110", "00111010001010110110", "11010101111011100101", "01001110000011110101", "11001001110010100111",
		 "00111110101011111101", "00111110110011001000", "10100001100011111000", "10110110000110000110", "01100110010011100100", "00110101111100101001", "11000110011100110111", "11011010000011000110", "01000101111011110111", "10111010010011111000", "00111010010100010111", "01000001100011100101", "01000101111011100101", "10111110100100110111", "01001101111100110101", "11000010111100101000", "10111110101100001011", "01111101110100111001", "01000110111100011000", "10110010110100101010", "00110001110011110101", "10110010000100000111", "00111010011011101001", "01011110011011001001", "01001001110011101010", "00110111011011000110", "11011101110100011010", "11000110001100010111", "01000001110100100111", "11000010110110101011", "10111110000100010110", "11001010111101001000", "01011110110101000111", "11110101111100110110", "00110001100011000110", "10111001100110001000", "11000001100100000111", "00110110010011000110", "00110001110100100111", "01010010111101110111", "00110101110011010110", "00111011000011011001", "11010010101011001000", "10110110101100000111", "01011110100100001100", "00110111011100011000", "00101001110010010101", "10110011000101111010", "01000001111100100011", "00101110100101011010",
		 "10110011110100010110", "00110110010011000111", "10110110000100001001", "01000010000011111001", "00110101110100101100", "01000001100110000111", "01010010000100011000", "01000010110101000111", "10110010011011100111", "01000010011100000110", "01001101111100001001", "11010101111011001011", "11000110000011110110", "10111010111011011000", "10110001101100100111", "00111110010011110110", "00111001110100001000", "00110110000100110110", "11001010001101110101", "10110110101100111000", "11011010000100010111", "01001010011100010110", "01010110001100110101", "00111101111110101010", "01000010001011101000", "10101010101011000111", "11000101110011101000", "00111110001101110101", "01001010011100101000", "11000110001101110110", "10101010011100001001", "10110010001100110111", "11000101110011001011", "10110110011101001010", "00110101100100000110", "01000001110101100110", "11000010011100011100", "10101110010101001000", "10110101110100101100", "11011110110100101001", "01001010001101100110", "11100010000100010101", "00100001001100000110", "00110010001011100111", "11010101111100001001", "10111010010101011000", "00111101110101000111", "10111110110100000111", "00111010001011110110", "10100010011100010111",
		 "10110110001100010111", "10111010011100001110", "01001110010100001001", "10101010001100101000", "01011010100100100110", "10110110000101110111", "01001110110100110110", "10101010101100101111", "00110110101100000100", "10111101100011001001", "00111010000011011010", "10101110100011101000", "11001010110101000110", "00111111000100001000", "10111101100110110110", "11010101110100001001", "11000001110100011101", "11000110001100111000", "10101101110011111000", "01000110101100010110", "01001001110011111010", "10110010010011110111", "01010010000011110101", "11101110100010100101", "01001011101011010111", "11000110011101001000", "10111110100101011000", "11000110001100001001", "00110010001011100111", "10110010001011001000", "01010010000101001000", "11000110000100111000", "11001110011011111010", "10111101111101101010", "10111010010101000101", "00111110001011011001", "01010110001100011000", "00110010100100000110", "01111010111011010110", "10110110000100101001", "11000101111011110111", "10110110001100001010", "10111110100100011000", "00111010001011100111", "00100001100010100101", "01001010011010111000", "10110010011011110111", "10110110100011100101", "01000001110101000101", "01000001110101100101",
		 "10111101101011000101", "01000010100100010100", "10110010001100111000", "00111001100011000101", "01001010011100010100", "00110001111011011011", "00111110000011101001", "00111111010100000111", "01000101010011111001", "10101101011011100111", "10111010000100101001", "10111110000100000111", "11001110010100010111", "01000001101011100111", "01101110010100001010", "11000110001011111000", "11000110001101110110", "00101001110010110110", "00101001100100100110", "00101001101011100111", "11011010001100001001", "00100010001100011000", "01000101100011110100", "00110001100100110110", "11001010011100011000", "00110101110011010111", "00111101110100111000", "11001010000100101010", "10111011010011100110", "01000010100100000110", "11000101110100000110", "01001010001011110101", "10110001110110010110", "00111011111100001001", "01011010001100110101", "11011101110110110100", "00111010000011001000", "01010001111100001000", "01001110000100010110", "10100010001100011001", "10111001111101000111", "01001010001011110101", "10110001000100000110", "01011011000100010111", "01101010010010110101", "01001001111100101000", "10111010001011000110", "10110110001100101101", "11000110001100000111", "00111101110100010101", 
		 "11000110001100101001", "01111110000100001000", "11000010010011101000", "01001110001101011001", "10111110000100101000", "10110101110100111100", "01000110010100010101", "01000110010100001001", "11001110010011111010", "00100110001101111010", "10110010010100111100", "01010110001100010110", "10111010101100011000", "11000111011100101000", "11001010011100010111", "01000010001101111100", "10110001111011100111", "01000110000011100111", "00110111101100110101", "01100010010100110101", "11000010011111010111", "01000110100100011001", "01001010101101110110", "11011010010100110101", "11011101110011101000", "11001010000100100101", "01001110000100011010", "11011110010100101010", "01001110001100011001", "10100110001101001000", "11001101110100011010", "01000111011010100110", "11010010010110011100", "01000001110101001001", "00111010110011101001", "00011010101100000110", "01010001100100000110", "01000110100101000110", "11000110011100100101", "01001110101101010111", "10111010101100101001", "11000110110100011000", "01001010010110011001", "10110110100100001011", "01000010011111011001", "01000011110011110110", "01011111010100010111", "01001110011100011001", "00101110000011001000", "10111010010100101000",
		 "11000010101100110111", "11000110011100001111", "11000010001100001000", "11000010101100000110", "11000010110100110101", "11011110001101110110", "00110110010011010110", "11000010100100000101", "00111001110101101001", "10111010100100101010", "10110001110011100101", "00110110101101000111", "11000001100100100100", "01000010011011111000", "01010001110110000101", "01000010010101010110", "00100001110101011010", "11010010000101000100", "01000101110100010111", "01000010000111101011", "11000010001101110101", "00110010011101000110", "01001110011100101001", "00111110110100111010", "01000010101101100101", "01100010001100101001", "00111110000111110110", "01001110011100110111", "11000110010100011000", "10111110011100110110", "10111110110100101001", "10111010100100111000", "00110011011111000111", "11011110001100010111", "10111110001100100110", "00111010001110010111", "11000010010101010100", "00111110000100000111", "11101110111011110110", "01001110010100011000", "10110001111101111001", "11001110010101111010", "01011010011100000111", "01010010110011010111", "11000010001100011101", "00111010001011000111", "01000010001100001000", "10111110000011100111", "10110101110011111010", "01000010100101010110",
		 "11000110000100000101", "11101110101110011001", "00110110101110000111", "00111010100100010110", "10110011010100001001", "00111010101101000111", "01001010001100000101", "00101010010100000110", "00111111100110110100", "01001010010010100111", "00111010101100010100", "11001010000101111000", "01001110001100110111", "01000010001100111000", "00111101111100011000", "01001010001100010110", "01010110111011100100", "01000110011100101010", "10101001111111001000", "10110110000111011000", "01011001111110101011", "11011010101101111000", "00100010010011100110", "00110010110100011010", "00111110101101110101", "11000110010100000110", "10110101111011101001", "11001101110101011000", "01011010110100110100", "00100111010101001011", "11001010011100010110", "01000111001100110101", "11011010011100011110", "01000111000100000110", "01000101101011011001", "00111010001110110111", "10110010101100101000", "11000110110100010100", "00110001111100100111", "11100010110100101011", "00111001010100010011", "00111001010100110101", "00101011001111000101", "01001001111100110111", "01000010011101011010", "00110110001100010111", "00111010010101000100", "01010110010110110110", "11001110000011110101", "11010110000100000110",
		 "00111110011011101010", "01000001110101001000", "10110110011011101001", "01000111011100001100", "01010110111101111000", "01000110001100100110", "11010110000101010111", "11000010001100100110", "11000001111011100110", "01000010000011100101", "01010110100100010101", "01011110011100110100", "01000001111100000101", "10110010011100010111", "01110010001100110101", "10111101110100101010", "11010110001100001000", "10100101111100001000", "10101110111100110101", "00110101110100100101", "11011101111100010110", "10100001110110011110", "00110101111110000100", "01010010000101011000", "11001101100100110111", "10111110101011111010", "11010110000010101000", "11000110001100001001", "01000010011011110110", "01000010011100111010", "01000110101100100110", "11100110010100111011", "10101110000100011001", "11000010001100000110", "00110010010100110100", "01000010000100011001", "01100110110100011001", "10101011011011110110", "10111101111101010110", "00111010000011110101", "11000010000011000110", "11010001110110000110", "11001001110101111011", "00111110111011110110", "11010110101100000110", "01001110001011110110", "10111010111100100101", "01010101110110001010", "11000010001101001010", "01001110110011110111",
		 "01000110001011111001", "01000110010100000101", "10110110001100000111", "11000110011100100101", "00101010011100011000", "01001010100100100100", "11001110011101111011", "11000010011100011001", "10101010101011001000", "01001010010011101001", "10110101110100111000", "00110010101011110101", "11010110100100110111", "01011110010100001001", "00110010100100010111", "01011110000011100111", "00110010001101001000", "00110001111011100101", "01010110000101010111", "11011010010101011011", "10111010000101001110", "01000001110101011001", "01000010011110100011", "00110110110100101000", "10111001110101001001", "10101001110100011000", "10100101101100001000", "00111101101110011000", "11010011111100000111", "01000010010110101100", "10110010101101110111", "01010110010101011001", "10111110010111111001", "10111010010100001010", "00110010000100010110", "10101001111100000110", "11000001111100101011", "10101010001101111000", "00111110010100100110", "00111110111101110100", "11000110101100000110", "01001010000101010110", "00111001011100101010", "11001110100100100111", "01100011110100011010", "01000010011101000111", "00111110011101000100", "10110110011100111001", "11011010110101111001", "00101110100100101000",
		 "01001110111100011010", "01010110010101011001", "01000011000100011000", "00101110011110010101", "10110101111100011000", "10110110000111111000", "11000010010100001101", "00111110011011100111", "00100011110100000100", "11101101111011110111", "01000001111101011011", "01001010011100111000", "10110110101100101101", "00111110000100000111", "00110101110100010101", "11000101110101110111", "00111010101100000101", "00110010010111110110", "10111110001101110111", "01000110000100010100", "10111010001101000101", "01001110011100110100", "00111101110011100111", "11011110000011110100", "10111110001100010100", "10111010001100001001", "11000010011101111001", "10111001110100001001", "01010110010100100101", "01010110010100110110", "01000010101100001000", "00110010000101110110", "01001110010101001010", "11010110000100111000", "10111110001100000111", "01001101111100111001", "01000010011100011000", "00111110000100001000", "10111110001100010110", "10110010011100000101", "01010010010100110111", "10100001111101011010", "01000010010100000110", "01110010111100010110", "11001110000011110111", "00101010010101100100", "01000110101100100111", "10110010100100100111", "01100110000011111000", "01000010010011010111",
		 "11001101111100110101", "01000110100101010101", "00111010100101101010", "10110101101011111101", "11010010011110010111", "10100010010100010111", "11011010010011000110", "10111110101100011000", "10111011101100001000", "10110101111111011001", "10110010100100001000", "11001110001011111000", "11001110010011110111", "10111110111101001010", "01010010101100101000", "11001001111011101001", "00111110010101000110", "11000010010011100111", "11001110000101011010", "00101001101101001000", "01000010110100001000", "10111010000100000110", "00111010010100010101", "01001010001100000111", "01001010111101000111", "11000110000100000111", "11000010011101011000", "11000011001100111001", "01000001110100010011", "01000110100100010011", "01000110011100000111", "10111011001100111011", "00101110011110000110", "01100111101011111011", "11001101111100011001", "01100110011101010110", "01001110011100110110", "01001110001100001010", "00111010000100010011", "11000010001101100110", "00111110011011010100", "00111010111100010101", "01000010011100000111", "01010010001101011000", "00111110100011000100", "10110010101101101011", "00101001110100110110", "11000110010100000111", "01000110000100110110", "00111001111011000110", 
		 "10111010101101001001", "00110101100100001100", "11000001011011111010", "11001101111011111010", "10111110110101011010", "10110110001100101000", "11010010000011110110", "10110010000100011000", "10111110100011110111", "01000010000100111010", "10011110101101100110", "11000010010100110111", "01111010001100010101", "00111010110110010111", "01001110101100100110", "11010010001011100101", "00101110000100110110", "00101010000011100110", "11001010000101010110", "01000111000011010011", "00111001111100110110", "00111010001100000111", "01001110001100110111", "10100010100100000100", "00111101110011100100", "10111001100100110110", "10111101110101110111", "11010010001101010101", "01000011011101100110", "01001101110110001001", "01011011101100111010", "01000011001100010101", "10110010010011110111", "00111001111101010101", "11000011000110000111", "10100110100011110101", "10110101101101010100", "01000010100101100100", "11001110000101000101", "10110110100100110110", "11011110000110011011", "10111101111100001001", "00111101011100000110", "01000011001100101001", "11010110001100111001", "00110110010100010111", "01001001110101010110", "01000010101100011000", "10111110011100101000", "00111010000100001010",
		 "11001110110100110111", "10111110111011001000", "01000001111011101010", "00111110010100010110", "01000010010100110111", "01000110001111000110", "10111110110011110101", "11100001011011100011", "00101011001101011000", "10101011110111110111", "10111110101101000100", "11001010100011100111", "01000001110011110100", "01000001111100111101", "01000011000011110110", "01000010101101010101", "10100101010100001001", "01000110001100010100", "00100010010011100111", "01001101111100001011", "00111010001011010111", "11001010011110110011", "10111010011100011000", "11000110100100101000", "11000110001100100111", "01110010111011110101", "01001110010100010111", "11000010011100111000", "01001010011100010101", "01000111001101101000", "10101110000101110111", "00111010111100001001", "10110110011011000111", "00111110011011011000", "01001001111100000100", "00110010011010100101", "11000111010011110110", "11000001111100000101", "10111110101100101001", "10110001110010100110", "10110001010101010110", "01010010101011100100", "11001110001011010111", "10111111000101110111", "01001101110011101010", "10101010010100001000", "01010010000011101010", "01000010000010100101", "01001110001011101000", "00101001110011010110",
		 "10111010000100100110", "01011001111110000111", "00101010011011000110", "10110110111011100100", "10111110001101001000", "00101110001011100100", "00110010000100010110", "00100110010011100100", "01011001110100010100", "10111010100011010101", "00111010011100000011", "01000110001100011000", "01000110011100000101", "11010110001011010111", "00111001100011011000", "01111110111101000011", "11101110011011100111", "10111110010100001011", "10101110010011101001", "10100111000100111000", "10110110101011010110", "00111010001011110100", "10101101111100011001", "11010010100100101001", "10101110111101110101", "00110110101011100101", "00101001011100111001", "11000101110101010101", "00110101110011100111", "10011101101011111001", "11001110100101110101", "01001001110011110100", "10110010001101010111", "10101110000100010110", "00110001011100000100", "10111101110100111001", "10101110011011101100", "10100010010011110011", "10101001010100101000", "00111010000101000110", "00110110010100000011", "10111101011011110101", "00110110011100000101", "00110010010100001000", "01010110011100110101", "01001001111011000011", "11001101101110000101", "01000001100111110110", "00111010000011000101", "00110110010100010110",
		 "01010110001100000101", "10110101110100001001", "10110010000100101000", "00011111001010100110", "00111010000011100101", "10110010111011100101", "11000010001101011000", "10101110111101000110", "00111110011011010110", "10110111010100010110", "01000001111101010111", "11010110011100000101", "10101101010100000101", "10111110101011101101", "00110010001011110010", "10101110000100011100", "11000110010011010111", "00110110101100111000", "00111010011011010100", "00110110010100110110", "10111001110011110110", "00110001010111001001", "10111001111101010011", "11000101111011111000", "10111101110100110110", "10011101111100011001", "00101101101011101011", "10101110000011010100", "10101101110100111000", "00110001110010100111", "01001110101101000100", "11000101100011000110", "11001001111101001000", "01000110011100010100", "00110110010100100100", "10110110011101001000", "11000110011100010110", "11000010000101100101", "10110101110100000100", "10111110000011110111", "00101010100011010100", "01000010011110110010", "10110101111011111000", "11001110011100110011", "11001110010011010100", "11001010011100010011", "11000110010011100110", "00110001110011001011", "00111101110100001000", "01000110001011011000",
		 "11000110000100001010", "10110010000100000101", "10111010001011101000", "00110101101100001000", "10111110011100010111", "10101001110011101000", "11010001110100010111", "00100110001100111001", "10100001110010000110", "00111010011011111000", "10101101111101000110", "10100101011011010110", "11000010000101110110", "00111010110100101000", "00110110000100001010", "01011110001100110011", "10111010000101110110", "00110110101100110011", "11010010001100010110", "11000010000101111000", "11001010011100101001", "11011001111011100101", "01001011110100010100", "00110101100100101000", "00111010010011010100", "00100010101011111000", "00100101100101101010", "10011001111011110111", "11000110000101101010", "00111010011100011000", "00101110010010101000", "11010110000011101001", "10100110010100111000", "11010010000101111010", "01111010000101010100", "01000010001100011000", "01000010001011001000", "10111010010101101001", "10101110110100010111", "01111110011100110110", "10101001111011010101", "01100111010100110111", "10110001111100110101", "01011011001010100101", "10111010100100101010", "01011001111100100100", "10101101111100100110", "00111110000011100111", "01001010001011100101", "00100101110100110110",
		 "10111010010100000111", "00110010010100011100", "10111101111100111001", "10100110010011100111", "00100001100011110111", "01000110011101110111", "11000010000011101000", "11010010000100011000", "00011101110110100110", "11000101011100000101", "11001110000100100110", "10111110011100110110", "11001010010010101000", "10101001110100101000", "10100110100100010101", "10110110000011101000", "00101001111011100110", "00110110011100111001", "10111110001100110111", "10101010101100100111", "10110110100100100110", "10101110011010110111", "10111101011011100110", "11001101100011000111", "00110010100101010101", "01000110000011111001", "11000110000100001000", "10101001101101001111", "00111110010100110111", "10110110100100100110", "01011010101100110110", "00110010000100001000", "10111010101100000110", "01111110100011110110", "11001010010111100110", "01010110001101111000", "00111010000100110110", "10110001111101000100", "00111001111100000110", "10011010001100001101", "10110101111100010110", "10011001111011111000", "00110010000101000101", "00101001110100000101", "10101001111100100011", "01001110111100000100", "11000101101011011001", "00101110111110000011", "01001001110100101001", "00110110010011101000",
		 "11000010011100000110", "10111010001100010101", "00110010011100011000", "10110101101100110110", "01000001111100010100", "11001001110100101000", "11001001111010001000", "01000010001101001000", "00111101101101011011", "10101110100100111001", "00101010001100000110", "10101110010100010110", "00111010001011111000", "10100010000011100110", "11000101111100111000", "00110001110101010010", "11010110010011110110", "10110010100011001000", "00101110101011101000", "00111010010011100110", "11010010000011111001", "00100010011011100111", "00110010000011110111", "00100001101100111011"); 
		weight_ROM(3) <= (
		 "11000010101100001000", "00111010100100101000", "01000001110100000111", "01000011001100001000", "01000001111011101001", "10110110101100100111", "00110010010100010101", "01100010111100001000", "00101010000100100111", "11000010000100101001", "00110010000011100111", "11000010011101001001", "11001001110100111001", "00111001111100101000", "01001110001100011000", "11000010011110011001", "11001010011100001000", "11001010010100011000", "11011010110100101100", "11001111001100011000", "01001010100111101001", "10111110001100001011", "01100010100100000111", "00101011001100100110", "01001101110100000110", "11010110111101010111", "11000010110100110101", "00110010001100110101", "00111010000100011000", "10111110000100101010", "01001010011100010110", "00111010000011000101", "10110101111100110110", "01001010011011111000", "11000111010100010111", "01001110010011110111", "01000010000100001000", "01001001110101010110", "00111010000101000101", "00110111010100000110", "00111101111011100111", "00111011011101000110", "01000110000100101010", "11000010100011101010", "01010110010100011000", "11000010010100101000", "00101010000100111001", "00111010100011110111", "00101001110011001010", "10110010001011101000",
		 "01001111101100011000", "01010010011101011000", "01000110001100010110", "00111010001011101000", "01110001110100111010", "01000101110100010111", "01001010110100000111", "01001111001110001011", "01000010000101111000", "11000010011100000111", "01010010100100111000", "01011010010100111000", "00111001110011100111", "10101010110100110111", "10110011111100111010", "01001010111100011000", "00110010011100101000", "00111110000101010110", "01010011000100000111", "01001010010101011001", "00111111011100011001", "01000110000100000101", "10111110010101110110", "10110001111011101010", "00111010000100101000", "00111010001100101000", "00111010000100010111", "10111010011100010111", "01001010100100011000", "00111110010101001001", "01000010101100101001", "01001110100111101011", "10101101100101001000", "00111010000100011000", "01000110100101110101", "01000110000011101000", "01011110101101000111", "11001010000011000111", "10111110000100110111", "11000010000100001000", "11000001111100101000", "11010110000011100111", "01011010001011100110", "11010110101100011001", "01001110101100111001", "01001010010100000111", "11000001110100111010", "01001010001101011001", "00111110100110110110", "11000010010101010110",
		 "00111010010101001001", "00111110000100001011", "00101010000100100111", "00110111010100101000", "10110101110011011100", "01001010000100011001", "11001011001100110111", "00101110110011100110", "00111010100100010100", "00111110100011100101", "11001010010011111000", "11001010000110010111", "01001110011100011000", "01001110010100111001", "11010010100100001000", "01001010001011110101", "01000111000100011001", "10111111001100101001", "11000110001101001000", "01010110011011001000", "11001110100011110111", "10111010011100101010", "01011010111100011001", "10110110101011101010", "00111010100011100110", "11101110011100010110", "00111110101101001000", "00111001111100100111", "01010011000100010111", "00110101101100000111", "00110110010100011000", "00111110001100101000", "00110001111101001001", "01010110000100110111", "11010011110100011001", "10101011111100001111", "10101110111101100111", "00111010100110111011", "10111111001111000111", "00111110110111101001", "01000101100011100111", "11001110111101110110", "00110110001101101000", "00111010101100000110", "01001110001100000111", "01001010011101011000", "01000110001011100110", "01001110011100100111", "00111111001101010111", "01000010000101000111",
		 "11001010010100001000", "00110010110100001000", "10110001110100000111", "10110111010100111001", "11000010010011100110", "11001101101010101000", "01010110010100110111", "10111001111011101001", "11010010110100111010", "11000010011101101000", "00111010111011100110", "01000010000100001000", "11011110100101000101", "11011010001100001001", "10101110010110110110", "10111110000100001000", "01001110111110011000", "11011010001100001011", "01011010001100001000", "01011010011011111001", "01001010001100010111", "10111010010100011001", "01000010000100001010", "01000010010100111001", "11001010001101101000", "11001010011101000110", "11001110011011101010", "10111010011100011001", "11001010000011011001", "11000110101100111000", "01000010001101010111", "00111110000110110110", "00111001110100111000", "01001010011100010101", "11001010100101000111", "00111110101101011100", "11000110010100000111", "10111010000100000110", "00110010000100100110", "11001010101100011001", "01000110011101111100", "01000110101101100111", "10110010000101001000", "10110101110100111000", "01001110100100010111", "01001010001100001000", "01000110000010101001", "11000110100100101000", "11001110011101100101", "01000110001101000111",
		 "11010011011110111001", "00111110111100001001", "11010110000100011001", "00110010000100001000", "00111101111011100110", "11010001110111110111", "01000010101100110111", "01000110000100001001", "10111110011110000110", "01000010001101001000", "11110110111101111000", "11000010011111011000", "11010110000011110101", "11000010011100110111", "01000010001100101000", "01000110011100110111", "11101001110101011010", "01010011101110100111", "11000010001011101001", "10110011011100111001", "11000110001101001000", "11010110011100010111", "11011010100101110111", "00111101011100011001", "01000110100100111001", "10111110000101000111", "10110101100011100111", "10111101110100110111", "00111010100100000111", "01101010011101011000", "10111110010100100111", "10110010011100001001", "10111110000011101011", "10101010101100001010", "01000110000100011000", "01001110101011100111", "10111010011100111100", "10101010010100001001", "11000101101101101001", "01000010000100110111", "01000011010100111000", "10111110100011111000", "00110010001011101000", "01001110101100001001", "11011110000100011001", "10111010000101111100", "01000010000100000110", "10110010101101101000", "00111001111100010110", "10111110001011110111",
		 "11001010111100011100", "01000010001100011010", "01000010001100001111", "11010011001101101000", "11001010011100100111", "11000110000100111010", "11011010010100101100", "11001011001110011000", "01000011001100101001", "01001001100100000110", "11000010000011110111", "00111010111100011001", "11000110001100101000", "11001010000011101000", "01000010000110101001", "10111111001100001001", "10111110010011100111", "00111110001101110111", "11001011001100111001", "00111010010011111001", "10111110010101011000", "10111010011110011000", "00110010100100110111", "01000010000011001000", "01001110001110100111", "01011110001100110110", "10111010111100001001", "10111110000101000111", "00111010010101111000", "11010110001011000110", "01011010011100101101", "11010110110101010111", "00111110000101011010", "11000010110101001000", "10111010000100001001", "00111111100101110110", "00111110000101011011", "01000010000101111001", "01001010101011110110", "00110010000011100111", "11001110011100001010", "01011110001110000111", "01001110000101011001", "01000010011011111000", "00101010010011100111", "01010010000110010110", "01011110100111001010", "01000111010101001000", "00111011001101001001", "11001111010100001001",
		 "01000010011100000101", "11001110010101011000", "01100110001110001001", "01001110000100000111", "01001010001100010111", "01000010011101001001", "01001010100011101100", "01000010011100001001", "10111101110101001000", "10111110000011111001", "10101010001100111000", "10111001111100001001", "01000110000100011001", "10111010101011101000", "00110011111101000111", "10111010101100010110", "10111011110011110101", "00111011110100010110", "00111010000101001000", "11001110000100011010", "00111010001101001000", "00110001111011111000", "11100110000100001000", "01001010000100011011", "11001011000101111000", "00111101110011110111", "11001110011101110110", "01001010011101011000", "11001010010100101001", "00111110100100011000", "01010110001100001010", "01111010101100101010", "10111010111011101011", "00111010011100000111", "01101110001100010101", "11001101100100011000", "00101001110100001001", "11000010000011111010", "01001010010011101000", "10110010011100011001", "01100010001101001000", "01000010100100110110", "11100001101101101000", "01000010110100001001", "01010111000011101101", "01001110101101011100", "10110010001100001000", "11000101101101011010", "01000010010100000101", "00111101110100010101", 
	 	 "11010011001100101001", "01001010100100001000", "01001010100100011010", "11000010000100001000", "00111110011100101010", "01001111011101011000", "11010010101100011001", "01000010000101011100", "11000010010101001010", "01010110011100011001", "11001110010100011011", "11000010011100110111", "01010010010100011010", "01010110100100111011", "11000101110100111001", "10111110001100001000", "11001111001100010111", "01000110010100001001", "01000101111101101000", "01001010000100101000", "01000010001100001001", "11000010000101001011", "01101010000101101000", "11000110010111011010", "11000010100101011001", "00111110010100100111", "11010110011100001000", "11101010010100011000", "11000010001101000111", "01010010111100111001", "11001010000100111000", "11001110100100011010", "11010101111100111001", "01000001111101001001", "11000110001101011000", "01001110011100111001", "11000110110011111010", "11010110110100011001", "01000011111110001000", "01001011001100001010", "11010010010101001011", "11000110010101011001", "00111110000100101001", "01000110010100011000", "01001010111101001011", "01010110011100011000", "01011110010101001011", "01101010110100101001", "11000001110101001001", "00111010000101001011",
		 "11011010000100011000", "11000110000100111011", "11100010010100101010", "01001110011100000111", "11000010011100110111", "10111010000100111010", "11011110011100101000", "11010110101100101001", "01001110001110001010", "11000011000100101000", "01011001110100111011", "01000010001100101000", "10111010100100101001", "01001110010101010111", "11001110001100111001", "11000011001110111000", "11000010001100011010", "11001010010100111001", "10111110101100111000", "01000010100100001010", "11011010100011101001", "01000110010100101010", "11000001111100000111", "01000010011100011101", "11001010010100011000", "11001010001100011010", "11011110001101001000", "11010010100100001000", "11000010000100101010", "01010110001100001000", "01010010111100011000", "01000010011100001111", "11000010000100011001", "01010111001100011001", "10111010011100011001", "11011011101101001000", "00111010111100101000", "10111110011011101011", "10111011000100111000", "11100110101100011010", "01001010101100011000", "11110110011101001000", "01101111100100101010", "11011010000110101000", "01011010101100101001", "01000110001101001000", "01010110011100101001", "11011110000100101001", "01000010110101101010", "11001010010100011000",
		 "01010010110100001000", "01000111001100001000", "01010001110100101100", "11001011001100011000", "11000110001100101000", "11010110001101001000", "11000010000101010111", "01000110000101011001", "11001010011101100111", "10111010001100011100", "11011010100100111010", "11001110000100101000", "01010010001101101000", "01101010010100111001", "11001010001100111001", "11000010010100111011", "01001110011101001001", "11000001110101011010", "01011010101100001000", "01001110110100011010", "11100001111110001010", "11011010110100111000", "01011010100100011000", "01001110011100111001", "01010110011100011010", "00111110001100011000", "01000110011110101000", "01000110101110111011", "11001010110101101001", "11000010000110111011", "01010110011100101001", "01000010101101100111", "11000010010100101001", "01001010101100001000", "11010010011100001000", "01011111010100101001", "01001101110100101001", "01001010011101001000", "01010110000101111100", "11001110011100001010", "01000010001101001001", "01100110011110111001", "11000110011101110111", "01010110100100111011", "11001110011101111001", "01001110000101101000", "01000010000101011000", "11010001111100101001", "01000010011101011101", "11100010000100101010",
		 "11110010110101111100", "11001001110101011011", "01000110010100111000", "11001110011101101001", "00111110101110100111", "11010010011100110111", "11010010110100111000", "01000010001100101000", "01000010011110101000", "11001110010100001001", "01001001110100111011", "11010001110110011010", "01001110100100000111", "01000010110100111000", "01001101110110111001", "11001010100100001100", "11010010001101001101", "01011110011100011011", "01001110110101000111", "00111110000100111000", "01001101110100111010", "11010010000101111000", "01010010100011111001", "00111110010101100111", "11001110000101001001", "01011101111100111001", "01011010010111100111", "11010110000110001000", "11001110100100001011", "01001110000100101001", "01010010000100010111", "11000010011100101111", "11010010001100001100", "11001101111110000111", "01000110001100101010", "01001110100101101100", "01101110010100101001", "01011110011100100111", "01011110010111101011", "01000010011100111000", "11000010011100111010", "11010010010111111010", "01000010000100011000", "11000110001100100111", "11010110111100101000", "10111010010100011000", "11010110010100101001", "10111010100100101000", "11001110010100111010", "11001110010100011001",
		 "01010010100100001101", "11001011010100010111", "11001010010111111011", "01000110001101001010", "01001011111101011000", "01010010000100001001", "01000010001100011001", "11100010001100001001", "01001010110101111001", "11011110000110101011", "01111110100100101000", "11000011001100001001", "00111011010100011001", "11010011000101001000", "01001011100100101011", "01010110010100011000", "11000010100101001111", "01010110000101101000", "01001010000100001001", "11011010001100011000", "11000110011110111010", "01010010111101101001", "11000010101110111001", "11001010110101000111", "11010110001100011000", "01001110011100111001", "01010110101110001001", "11000011110100001010", "01001110000100011010", "01001110011101011001", "11011010111100010111", "01010110011101001000", "01010010101100100111", "01001110101011101011", "01100110100100001000", "01000010011110011000", "01010110010110001000", "11000001111100001000", "11001111000100111011", "01110110010101011000", "01001110001100111011", "10111110001101001010", "01010010001101101111", "01001010001100001001", "11001010010011111001", "10111010100101001001", "01011110000101110111", "11010001110011111010", "11000110010100001001", "01110111101110001001",
		 "11010110101111000111", "11001010000100001010", "11011010000100011101", "10111001110100000111", "11001110011100111001", "01000110011100011001", "11001010010101101001", "11001010010100001001", "10111011001100001010", "11000110101100111001", "01001010101100001000", "01000010100111101000", "01001101111110011010", "11001101110100111001", "01001010000100001000", "01001110001011101000", "00111011010100011001", "11011010101100111001", "10111010010101001000", "11001110000100001000", "01001010101101001010", "11011001110101011000", "00111010011100101001", "11000010101101001010", "01000010100100111000", "11010101111100111001", "01010110011100011000", "00111110110101011001", "01000101111100011001", "01000010111111001000", "11010110000100111010", "11001110011110101001", "11010010111100010111", "00111010101100111001", "11110010011101001000", "01001010000101001010", "01001010101100001000", "01011010000111100111", "11001110000100111011", "01000110011100000111", "01111110000100001011", "01000110111100111010", "11010010010111101001", "01000101110100011000", "11001110100100011000", "11010010000100110111", "11000110011101001010", "11011010010100011001", "01001110101100101000", "11001110001100101001",
		 "01000110010100011001", "11001110000100011001", "00111010001101011001", "01010110011110111001", "11001110001101001010", "11001010000101011011", "10111110010100111000", "11001110100100111010", "11011010100100111001", "11101010101100101001", "01000101111100011000", "11011001111100110111", "11011011000100001000", "11001010001100111101", "01001110000100101101", "11010010011100111011", "01011101111101100111", "11010010010100101000", "01101110010100110111", "11000101110101001001", "01011010001100010111", "01011010011100111000", "11000010011100011010", "01011010000100111001", "01001010000101001000", "11000111100101001000", "11100110000100001001", "10111110000101010111", "11001110101100101000", "01010010001100101011", "01010010000101001000", "00111010101011101001", "11000110001100111011", "01000110101100101000", "01000110010100101000", "11001110001100101001", "11001010100101011010", "11001110010011111011", "11010110100100000111", "01000010000100000111", "01000111001011110111", "01000110000100111001", "11000110001110011010", "11101110000101010111", "11001111001110001000", "01001110010100111010", "01001010101110011000", "11000110111100111011", "11001010010100001010", "00101010001011101000", 
		 "10110010101100101001", "01010010110100001110", "10111110101100011000", "11001110001100111010", "01111110111101011011", "11000110001100101001", "11000110001101110110", "01010010000100001001", "01000110100100011000", "10111110000100101000", "00101011000100011010", "01010110111011100101", "01001010010101101000", "11001010001100101000", "11010110001100001010", "01000011101100000110", "11010110001101110110", "11001010001011111000", "01001110101100101000", "01101110001100101010", "01010010010100010111", "11000010100100011001", "11000110011011111011", "01000110101111011010", "10111110011011100110", "11000010100100110100", "11010110010100011001", "11000010101101011000", "10111010011110101000", "10111010001100111010", "11001010101011101011", "11100110001011110110", "10111110101100000111", "00111010101100011001", "01001010010100110110", "11000110110011010111", "01000010000100101000", "00111011111100101011", "01001110011101000101", "01001010011100100110", "11010001111011111001", "00111110101100101011", "01010110001101001000", "00101010011100000111", "11001110010111101011", "00111110010011111000", "11101110000110001001", "01001101110101111001", "00110111000011001000", "11001110001100111010",
		 "01000110001100111001", "11100110110011101010", "01001010000100001000", "01001010001011101100", "01101010011110010101", "01000110010011000111", "01000110011100000110", "11001110010101000100", "11001010000100111000", "01001010010100011000", "01000010000101000101", "10111110011100011000", "11000110010100010101", "11000001110101011011", "01000111010100000111", "01001110011100111000", "11010001111100101000", "10111110001100100111", "10111110000100101001", "00111101111011101001", "01010110100011111000", "01010110010101010101", "01111101111111010111", "00111010101101001001", "01001010001100111001", "01001010000101101101", "11000110010100011001", "11000110001101101011", "11001010011100001011", "10111110010100010111", "11000010011100111000", "11000010001100101000", "01011001111110001001", "11011010011100000111", "01000010100011110110", "01100110000101101011", "11001110111101111000", "01000010000101100111", "10111010001100011000", "01000110001100101001", "01001110110110001000", "01001010111101000100", "01100010111100011000", "11001111001101010110", "01010010010111101000", "01010010010101110111", "10111111001101011010", "11001010101100100110", "11010110011110111100", "01000001110101011001",
		 "10110001110101001000", "11001010000100000111", "11000111011100111110", "00111010000100000111", "10110010010101001100", "11001101110100101010", "11001110011100111100", "01001110100101100101", "01001010011101011000", "01001111010100010111", "01001110100011011001", "01001010010101101111", "01000110001011101000", "01000110000111011011", "01000110011100101001", "11001010011100001000", "01010011000101111010", "10110010001100001000", "00110110010011111011", "00111010000101011010", "01001010100101001000", "11000010000100101010", "11010010101100011000", "00111101111011100110", "11100110011100000110", "01001010111100100111", "00110110010100101000", "01001010110100011000", "11000101110011110111", "01000101011100101011", "00111101111100100110", "11001110000100110111", "11001110101101111001", "10101110000100110110", "01001110001011100110", "11000101111100111001", "00111010000011100110", "11010001111011110110", "11100010010100111001", "01000001110100101001", "11110110010100101000", "01010010001100010111", "11000111001011100110", "01000010110100011011", "01001110111100101001", "01100110101100001001", "01001101110100110111", "01110010111100010101", "11011110010101000111", "10111110111100111001",
		 "11000110010100101000", "01000010010011000110", "10110111010100111011", "10111110011011111001", "11011110111100001000", "11011110010100100101", "00111010101101111000", "10111101111100101001", "01010011011011111001", "11000010011101100110", "01001010011100010110", "01011011000100100101", "10111110010101101000", "01001110001011101000", "01000110000100010100", "11000101110101111000", "11010010011100100111", "01000101100100111000", "00111101110100010111", "11000010011101110101", "01000110000100010111", "10110110101101011010", "01000110000011110111", "11101001110101001001", "01000010001100001010", "10111010011100101010", "01011010011011001000", "00111010101110111001", "01001110011010101000", "10110010011010110111", "01011010011100010110", "10111010010100110110", "00111010001100011001", "01000010110100110110", "11010110011100100110", "10111001110100001001", "01000110011011101110", "11000010010100111100", "01001010111100001001", "01100010100100011000", "00110101110110000101", "11010110010100010110", "11000010010100011000", "10111010110100101100", "01001010001100111000", "00111011111100010101", "01001010001100000111", "00110110000011000111", "01000010010100101001", "01000010010100001100",
		 "11001010010101101010", "11011110011100000111", "11000110001100111000", "01100110001100000111", "01000010100100110111", "11000110000011100110", "11011001110100011001", "00110110000100001000", "10110110101100111100", "11000010111101111001", "11011110000100111000", "10101010111101111001", "01011110100100101100", "11100110101100011001", "00111010001100111100", "01000110001101110111", "11000110000100011000", "00111110100100110111", "11000010000100011001", "11000010010101101010", "11000010000110111001", "11000110110100010110", "01000110110100010101", "11000101111110001001", "01000110001100001000", "01100010011101011010", "11010010100100001000", "10101110101101001000", "01010110000011101000", "10111110011100101001", "10110010001100101000", "11001110100100111001", "10111010011100011001", "10101010011011101000", "11000110010100010111", "11001010011011100111", "10101110100011111010", "00111010101100101000", "11010011010100011011", "01000011001100111000", "00111010010100111000", "01001011111100110111", "00110010001100110110", "11011010111011101001", "11101111001011101010", "11110010100101011000", "11001110011110111000", "11000010010011111011", "01010110010011111000", "11010110101100010111",
		 "11000010001011101010", "11000110001101101001", "00111010011100011001", "01100010010101000111", "01011110001101001000", "01000110000101000110", "01000010101011101000", "11001010001100000111", "01011010101101011010", "00110010010101011000", "11001010001100101001", "11001001110101111010", "11001110110100001001", "00111110011101011011", "11100011110101011011", "10111010011100101110", "01001001111101111100", "11001010011011101010", "01000110100100110111", "01000110000101011101", "11000010001100001001", "10111111010011100101", "00110010001101011000", "11001110000100011100", "01010101110100110110", "11000110000100110111", "01101110011100011000", "11000010010100010111", "00111110000100100111", "11001110010110010110", "11000110101100111100", "00110110001111000110", "11001001110101000111", "11001010011011111010", "11011010011100011011", "10111111001100111101", "11001010011100101000", "01011110001100001000", "11001010010101100111", "10101010100011111001", "11000010001101001001", "01001010101100111100", "01001010001111001001", "11101010010100100101", "10110010010100011010", "01010010000110010110", "01000010001101101001", "01000010101011101011", "01010010100011101100", "11101110101011101001",
		 "11010010010101100111", "11000010000110010111", "11001010111100101011", "10110110010100100101", "01110010010011111000", "10111110100100001011", "11001010010011101000", "10111010111101001100", "11001110101101001000", "11000101110101011100", "10110110011101101000", "10110010011101001010", "10111010001101011011", "01000110010100011010", "00111110001110011010", "00110010000101001000", "10111010011100011001", "10111110000100001111", "01000010000100000111", "10111011110110010111", "01010110010101001001", "11000101110100111000", "10101010011100110101", "00110110101100000111"); 
		weight_ROM(4) <= (
		 "10111010100100001001", "10111101111011101001", "11000001100100011010", "11001001110100100111", "11110011110100010111", "00110010011100000110", "10110001110011100100", "00110110000101001001", "00101010000100001110", "10110010010101001001", "10101010011101000111", "01011010000100010101", "00110001100101100111", "01011011010100011000", "11010010010100100110", "01001011000100111001", "10101110011100010110", "00111110001101110011", "01010010011101100101", "11001110100011010100", "01001010011100110101", "00101101110101000111", "01001010100100101001", "01000110001100011010", "11001101010011110100", "01001110001100010101", "01000010011100010101", "11000010000100010111", "01000010011011110011", "10100110011011101010", "10111010010100100111", "01000010100011110110", "11000101111100100101", "11011101111011110100", "10110010000011001000", "00100011011100110110", "10101010110100100110", "11011010011011110111", "00110001111100100100", "01000010010100111000", "10101001110100101010", "11001110000101000111", "00110101111111000111", "00100010001101111000", "01000001110100111011", "10101110010100100101", "01000010001011110100", "01011110000101011011", "00011010000011000111", "11000110101100001000",
		 "01001110000101111000", "10111110110110010111", "10111001111100100100", "11001110101011110111", "01000010011100010101", "01001010000100010100", "00111110100011100110", "00111010101101010101", "01001110110100110101", "10110110100011100111", "00111010000100110011", "00111010110100010101", "01001001110011110101", "00101010100101011001", "01000101111101001010", "01001101110100010110", "01000001101101111001", "10101010110100010101", "00110110001101101010", "10110110100100011000", "11001101110110110111", "00110001110011100011", "11000111000100011010", "10111110110100001000", "10101111000100010100", "00110110001011111001", "10111001111100010101", "10111010111100101010", "10111110010100011101", "10111110111101101000", "10110110010100001000", "11001110110101111001", "01000110011100101010", "01010110000011011000", "11001010100100000110", "11010011111011000110", "01000110100100100101", "01011111000100000101", "11000011001100100101", "10101001110010110111", "10101110101011000111", "11101110001100001000", "10111110001011111000", "10111011101110110100", "00111110010100100101", "10101010000011010111", "10100010100100010110", "11001101111010110101", "01000110000110000111", "11001010010100000100",
		 "01000110010100000100", "01000110010011100100", "01000001110011111100", "01000011001011110011", "10110110101100111001", "10110101110101010101", "11101110110100010110", "01100110000011010101", "11000110101100110100", "01000110100011000011", "11010010011100100010", "01001111011100111000", "01001110000100010111", "10110110001101101001", "01010110100100111000", "00111111011011011000", "10110001100100100101", "10110010000100011001", "00111111000100011001", "00110101110100001001", "01000110011101101101", "00110110011011000101", "10110001111100010111", "10111101110100011000", "10111101111110000100", "11000111001011000101", "00011110001100000101", "11001101101100101001", "00110110011100000101", "10111111001100011001", "10110110101100001000", "11010110010011010111", "00101101111100001001", "10110110000100000111", "10101001100100010111", "10110110000011101010", "10110010000011011000", "00100010101101100110", "00101001111110111010", "11010110010101001010", "00111101110110000110", "10101001001101000100", "00110101111011100101", "00110110010100101010", "11001110000101010101", "00110010101100010110", "00101001110011010110", "11010101110101011000", "11011010000100010101", "00111010001100010110",
		 "11010010001100010110", "01001001110011100110", "00110010010100001100", "00110110000100100110", "01000111000011100110", "10110110001010110100", "01010101111101010110", "00101001110100000110", "10111101111100011000", "00110010000011100110", "01100010001100010100", "01001010011100000101", "01000001101100001000", "11001011000101011001", "01000101100101110101", "10101010010100101001", "00111110010100001011", "10101101000010111001", "11000010111100010111", "10111010000101000101", "11000110101101010110", "10110110100100001000", "01111010001011101000", "00111011010101111001", "11000010101100011000", "10110001101100001101", "10100101111100111001", "10110110011100001001", "01100011010011100110", "00011110100010100111", "01001010010110000110", "11000101110011001000", "10101110011100011001", "01000110011100110110", "11000010010011101001", "01011010001101111001", "11000001101011111001", "00111110000011111001", "00110010011101100101", "11000010101100110101", "00111010010011100111", "00111110000110000100", "00110101101011110110", "11001010101011110100", "10110010001100010101", "00111110101101010100", "10110110010010110110", "01000110001011111000", "10111110100111000101", "10111110001100001000",
		 "01001110000100100110", "11001010010101000111", "10110110010100001000", "00111110110100010101", "11010101111100010111", "01001010100101000101", "11000010001101110110", "00110110000101011000", "10101001110100001000", "10101110000100011100", "00011001010011101001", "10111010010100010101", "10111010011011110111", "01001101110100001001", "01000001100100101010", "11011010000100010101", "10101010000100011010", "01000110100011101000", "11000011111011100111", "11001110010101011010", "00110011110100011001", "01000110101101010101", "11001010010100010011", "00100010001011100110", "10110111101101010101", "10101111101100001000", "10101111101100111000", "00011010001100000110", "11000110010100101000", "11000110001100011000", "10110001111011001001", "01001010001101001100", "10101110000011111001", "11000110010101001110", "10111101010011111000", "01010010011100010101", "00101010100011001000", "10101001111100101000", "00111111001011111000", "01100110101110000110", "00110001101100000110", "11000010000100111000", "00101001011011100100", "11001010100100111000", "11001110010100001000", "11000010000101010100", "10110101110101110111", "10110010111100001011", "11001010001101000111", "01000010001011100110",
		 "11001011000100001000", "10101010000100011001", "10111001111100101000", "00111010001101011000", "10110110001100001000", "11001011111101001000", "01010110101101001010", "11101010011100001010", "00011110001100001101", "10110101011100001010", "01000001100100100111", "11000110100101010110", "00111110110011000110", "00111010000100010111", "10110101010101110100", "11001101100100111000", "00101110011100100100", "00110101110100110101", "10110110001101000110", "01010010101101010100", "00110110001101000110", "01000110000110010110", "01010101101100101000", "10111101010011100111", "11000010101101010110", "10100110000100101000", "01001110001100111001", "10110110011100001000", "11000010111100000110", "10110110111100011010", "11001010010111101000", "10111001111100110111", "01010001111101010100", "01011010010101011011", "10100110000100001000", "01000010101100111000", "01010110010101110111", "00110001110100000101", "01000110000100010110", "10111001110011100101", "01000010010100011010", "10011010001100111010", "10110001111100000110", "11001010110100000101", "00100001110100100110", "10101110010110000101", "11001010010101101111", "00111111001100000110", "11010010000100001010", "10111010001100100100",
		 "01010001111100000101", "11001010100101010111", "00101010010101000111", "00110110010011100100", "00110110011110010101", "10111101111011010111", "11000110001011100101", "00110010010100100111", "10111010011011100110", "10101101110100001001", "10101110011100001010", "10101101111101100110", "11001101110100111010", "10100001101100001000", "10111001110100001000", "00101010000100000101", "01010001110011110111", "00101010110011100101", "00101001010100001010", "10110001101100000111", "01000010011101111010", "00101010011011001010", "00111010100100010110", "00111001110101100101", "10110010101100100101", "01000011010100010011", "00110001110011111000", "10111110000101000110", "00101001011110010110", "11010110000100000110", "10110010100100001000", "11000010010100101010", "00100001100111100110", "11000010010101000111", "11001010010100100111", "01000110001011110011", "10101110010101111000", "01010010101100111001", "10110010110101010101", "00110010100011111001", "10110111000011111001", "00111010100100100110", "00101110010100000111", "01000010001100011001", "11001010010011000110", "10101110010100010111", "00011110011011100110", "10101101111100100111", "00101010000100110100", "00111101110100010101", 
		 "01001010001101001111", "01000110001100000111", "01011010010100111011", "00110001111011110111", "10110010001011111010", "10100010111100000111", "11010010010011110011", "10110110010011111100", "00101010000100011001", "01000101111100100110", "01001001101100101000", "01000110100100101001", "11000110000100001000", "01000001111100010111", "00111110011010110110", "10111010000101010101", "00110010001011110111", "01000010110011111101", "00110001111100110101", "00111010000010111000", "11001010001011010111", "10110110011011110110", "01011110100100010111", "00111001101011100101", "00111101110011100110", "10111010101111000110", "10111110010101010101", "00110010001101010110", "00111010010101110110", "10101101110100001001", "01001110000100010111", "00111010000010000101", "10110101100100010101", "11010010011100010110", "10110101110100010111", "10111010000100011010", "01000010001101010101", "01011001111101001010", "00111010011011100100", "00111010000100000110", "00110110101011001001", "00111110011100011001", "01000001111011000101", "10101001111100011000", "01011010100100110111", "10101001110101000101", "00110010011011111001", "01000010000011110110", "00110010000100011001", "10101010100011101001",
		 "01000010011011110110", "01000110001100101011", "00111010101010101001", "11000001101100010110", "11001001111110010110", "00110101110011110110", "00111010000100010110", "10111010000100000111", "00110001111010111000", "10111001011011101000", "11000010001110110110", "01000001110111111000", "11001001111101000110", "10101101111011101011", "01000110111100001001", "10111011000100110111", "00101001000100000110", "01001001110100000111", "01010110001100001001", "01011101111100101000", "01001110001100110111", "00111101111100010110", "10111110100101010101", "10100110000100001000", "11000010000011111001", "11011110111100011010", "10110010101011001000", "11000110000100011000", "01010010010011010111", "01000010001011000111", "01000010011011100111", "11001101110100001001", "11001101011010100111", "11001110100101010110", "11000001111011101000", "11001001111011111000", "10110001110011110101", "11001110000011110111", "10111010001101110111", "10111010010011101000", "00101001111100110101", "01001001101101000101", "10111110011100000101", "01001110001100110101", "01000010000100011001", "00111001101011000111", "10101001101100000110", "01010001110011011001", "00111010001100010110", "11000010100100010100",
		 "01000010000011100101", "00111110010100010110", "00110010011101011010", "10111010000011100101", "10110101100011111001", "00111110101011001000", "11011010010101110111", "00110001110100000101", "00101010010100010111", "00110110100011100100", "00111010100100011001", "01010110010100110100", "00111010110101001010", "01000110001011100111", "10110110001101001001", "00111001111011100101", "01010010011011110111", "10101010110011001010", "01000101111011100111", "00110001111100001000", "11000001111011110111", "01001001101101110101", "11000101111100001011", "10110010011100001011", "00101010000011010101", "00111110010101000110", "01000111011011000101", "00110101010011110110", "00101010010011110101", "00110010001100101000", "01000010010101110111", "00111010100011010101", "00101001111101111000", "01000110010011110110", "10111101100100100111", "10110010000011101001", "10101010001011000111", "01001001101011101000", "00110101111110100111", "01011110101100010101", "00111110010011111001", "00110001101011010111", "00101001010011100101", "01000111001011000111", "01000110011011011001", "00111010100011110101", "00110110011011110110", "00101110011011100100", "00110010001101110101", "11000001110011000100",
		 "11001110101100011000", "00101010000010100101", "10100001110011000111", "10101001111011000100", "10111110000100110110", "10111101111101001000", "11011110100110110110", "10110001110011111011", "00110101111100011000", "00110010000011110101", "01000001111011100110", "00110001110011100111", "00100101111011100100", "11000110000101111001", "11000101111011110100", "10101110001100111100", "10101001100100111001", "10111111100100011010", "00101011001010110111", "10111101110100010110", "00110001100011010110", "00111010001100111001", "01001111101011001111", "11010010001011111000", "01000111000011101000", "01010101111011100111", "10111101100100011011", "10110101111101110110", "00110001110011000111", "11000010110011000101", "11000010111101001000", "10111101100100001011", "01000011000101011001", "01000101111011100111", "00110001110100010111", "10101001111011111001", "00111010001110100110", "00111010000011001000", "00110001110100000110", "11010101101101010110", "00111110000011110101", "00110110010011100110", "10111110001100011001", "10110111101010100111", "01001001111100100110", "11010010111011101000", "00110011000011010110", "10101010101011101101", "01000110000100100101", "00110110011100010110",
		 "10111101111101010110", "11001010010011100110", "10110110000111101010", "00111010010011100101", "00110101110100110111", "01101001101100110111", "00110010101100110111", "00111101110100011010", "11000110011011001001", "01000010001011100111", "01001101110100101010", "01001110001011101000", "11000010001100110100", "10111101111011110111", "10110010001011101110", "01010101110010101001", "00101001100010100111", "01000110100011110111", "00110010011100011001", "11010110111011010111", "10111010101100010111", "01010010011100000111", "11011110000100110100", "11000101100100101000", "01000010001010101000", "10101011001100001000", "10111101100011101001", "10111110011011110101", "11000001111101101000", "11000101111100110110", "10110010001011100111", "11000001100110011000", "10101110010011111000", "10101110100100101110", "00110010000011000111", "01000001110100000101", "10110110111011100111", "10100101110100101101", "10111101101101011011", "01000001110101101000", "00110001101011010111", "10111001111100010110", "00101010011100000110", "00110010000011101000", "10110010100100101001", "10111110000100000110", "00110101110010100111", "11000110000100111101", "00110010001100010110", "10101111001100011000",
		 "10100110011100001111", "01001010101011000111", "00111110101100000111", "11000001101100100110", "00111110000011100111", "10111110000101000111", "01111101110100101000", "10111101111100101010", "00111010101100000101", "10101101010011100111", "01001001110100011000", "01000011011011100100", "11010001111100000111", "10111010010101001011", "11010010110011010110", "11001001111110000111", "10110110100101011000", "11010110110011110110", "10111110000100011000", "00110010110011000110", "10111010001100110110", "10110010001100010110", "00110101111011011101", "00111101110011100110", "11000010000100110101", "10111110010011100101", "10111110001100011000", "11000101111100010111", "00101010001100000110", "01101110001100010110", "00111110011100010111", "01010101111011110110", "01000110111101101001", "10111010000101011000", "10110010000100000101", "01101010100101010111", "00111010000100110111", "00110001110100100110", "01010110011011100110", "01001110100011011000", "10111011001101011100", "10111110011011011001", "11001010100100101001", "00111010001010110110", "00101010000011100101", "10110110001011110110", "10111110101100011000", "10111110100011100111", "00111010001100101001", "10110001110101000110",
		 "11001101111011100101", "00111010011011110010", "10110010100101010111", "11001101100011000111", "01100001111100010111", "00110001101011000110", "00111110100011000111", "10111010111101111000", "01111101011011001011", "10101110001011011010", "10111101111101000110", "11000110100011000110", "11001101110011101011", "10111001100111100110", "11000110010011100111", "10111110001011010111", "11000110000011110111", "00111001100100110110", "00111110001011000111", "00101001011100000101", "00111010000110011100", "01000010001100000110", "01000101110011010101", "10111011001100110101", "01010110001101001000", "00111110000110110101", "10110110000100010101", "11000110010100010111", "10110110000011100110", "00111010000011101000", "00110110000101000110", "01001110010110010110", "10101001110011111000", "01010001111100011000", "00111010000011010101", "01001101110100110110", "01101001110010100101", "01001010010101001001", "01001010000110110101", "10110110011100001011", "00110010011011100111", "00111010111011010100", "10111010010010100101", "01010010011011111001", "11010110000011110111", "10111011001100011001", "10110010000100011001", "10110110011100010111", "00111110001101011001", "00011110010100010110", 
		 "10111101110011110111", "11000101110100001000", "10101001111010110111", "01001010100100011011", "10111110010100001000", "10101101111100101111", "01000110010101000110", "00101110011100010111", "11000010010101001000", "11001010000110111101", "10110010010011111000", "11010110010100100101", "00100001111011000100", "00111110001100000110", "01110010010100000100", "01000010001100010111", "01000110001100000111", "01100001111101010101", "00110001110101010101", "00110110010011110101", "11010010101100001111", "10011001101011111000", "01000110111100110110", "00111110110100000111", "11100101100011000111", "00110010001101000101", "11100110111100010100", "10111001100100101111", "10110110110100110101", "10110110010100001011", "11001110011100110110", "00111001101011110101", "01000101110100110101", "00111001111011010100", "11000101111100001011", "10100010010100011001", "00111001110100110110", "10101010100011100011", "10111001110110100100", "11100010011101100100", "10101001110100000111", "11000110010101101000", "10110010011100001001", "00111110010100100101", "11001110101101001000", "10110001111100010101", "01011111011101100100", "01010010000101000110", "00100001100100100111", "10111010010111101000",
		 "01000110001011100111", "10111101110101001010", "01000110000111100101", "10110110001100100110", "00111011011100000110", "01000010010100001011", "11011010001100110100", "10101010000100100110", "01001010101101001000", "10111001101011111001", "00111110100100110101", "00111010000110111000", "01000010000100010011", "00111001110100001000", "00111110010100110110", "11000110010100010100", "10111101110100000111", "11001101110100010101", "10110010010100000111", "10110111000011111000", "11110010001100001000", "00111110001011110101", "11001110011100000111", "10101001110100111011", "10101110000111110110", "11001111011100011001", "01010110000100110111", "01001010011011110110", "01000010101100101000", "01000010011100111000", "10111110011100000111", "11000110100100011000", "00101101110010101000", "01010111010100111011", "10111110110100000100", "00110010001100000110", "10111101110011100100", "00111110000100100110", "01000110010101010110", "00101001110011111011", "10101101110101010110", "10101110001110000110", "11000101100101100111", "10111010011100110110", "01001010001100101001", "01000010000011100101", "11100110001101100111", "10111010001011000101", "10101110011011101000", "00110001111100100111",
		 "10111010101100010110", "00110010010100000101", "10110001101100000110", "10110010011100110110", "00110010001100110111", "01000010001101100111", "00111010011100011000", "10111110110100101101", "11001010011110100110", "01000001111100010111", "01000110001100000111", "11011010000101010111", "01000110000100011000", "11000110111100101000", "10111001110100101011", "00111010011011111001", "11100010011100110101", "10110010011011101010", "00101010010100010110", "00110101100011101010", "00111110000011101100", "01011001111101000100", "00111110001100000110", "00111010011100001000", "01010011010011111000", "11010010100101110101", "11000110001100001001", "11010001111110010111", "10110001111011101001", "00110101111100011010", "01000110000100110101", "01001010101110000111", "11001110001011111000", "11001010100100010111", "10111001101100011001", "00101001010100011010", "10111101110011111001", "10110010010100000101", "10111010001100010111", "11101101111101100101", "10101001111100100100", "00110010001101000101", "10111001111101000011", "10110010100011111001", "01010111001101010110", "11000110000100110101", "00101101100010010110", "00110010001100010100", "01000011000100110101", "10101101111110100101",
		 "01010110010110011000", "00111001010011100110", "10110001111101011101", "00101110011101101001", "01000110011101011101", "01001001110011100111", "11011001111100010110", "01000011001100100110", "11000101111100011000", "00100110110011001001", "01000010110100110011", "01000110000011100111", "00100010101110010100", "11011010101101101010", "00111010110100010011", "11000010000100101000", "10101110101101111011", "01001110011011011010", "00110001111100100100", "10101101110101010111", "00111110010101010100", "10111101100100001000", "01000110000101011001", "11010110000100001000", "11001101111011110111", "00100010001100001010", "10101110100011011010", "01000010010011110110", "00111011000011000110", "00101010001011010110", "10110010001100100110", "11000110000100110110", "10111111010100001001", "01000010001100110101", "00110110001100100010", "00111010101011110111", "11000010101100001001", "10101110000100110101", "10101101011101001111", "11001110011100010100", "00110110100101100101", "01000010000110100101", "10111101101101001000", "10111110000101000101", "00110101111011100101", "10101110011100010111", "11000110010010100011", "11010110000100010111", "10110110101100100111", "11000101111011000110",
		 "11011101111101111000", "01001110000100000100", "01000110100110111010", "00110110011100000100", "10111110101101010100", "11000001110100000100", "11001010000100110111", "00110010011100110110", "10101001110100111110", "00111001111011101001", "00101001100100001010", "00110110000011010110", "11010010011100110111", "11011010100100101001", "10101010001011101000", "01000110010100000101", "01000110111100101000", "00110010111100110100", "11001010001100000111", "11001111001100101011", "01000010101100111001", "10111010100101100110", "01010110011110110100", "00110110000011101010", "01000001110101110100", "10100110010100000111", "00100101100101001010", "10111101010111010111", "11010110001100010111", "11011110010101000111", "00110101110011111000", "11000010000101000111", "10110101100011111001", "10110101111100111000", "00101001100100110111", "10110110101100110100", "10101001100100001100", "00011010010011011010", "10111010000101110111", "00111010010100100101", "01001010011110100100", "11000010010100010111", "11000001111100100111", "11010010000100010111", "11001011100100011010", "11000001111011101000", "00110001111011110101", "00110010100101001010", "01100001101101100110", "00101110001100001000",
		 "11001011111100101000", "10100101100100101001", "01000010001100101000", "00100010011100101000", "01100001100101000110", "10110001110100010111", "11001010000100111001", "01001101111100111000", "10101101100101010101", "00110101110011001001", "01000001111100111011", "11000110101100001000", "10111010011100000110", "10110010000110101001", "01111101010100010110", "01010110001100111001", "00101010001101010111", "10110010000100100111", "01010010010100010110", "11001110001101010011", "00111110010100110100", "00101101111100010111", "10111010001100000110", "01000001110011100101", "01001010001100110101", "00111110001100001000", "01001110100101011100", "00111001100101100110", "11101001111101010101", "00101010101011100101", "11000010101100110111", "10110110000101010101", "10111010011011111000", "11000110100100001100", "10110101111011100110", "11000110000101001001", "00111010010100101001", "00110101110101010101", "11001010001100001000", "10111010010011100101", "11001010011101001001", "00101011000100110111", "01010010011100110111", "00110010000100110111", "10101110111100010101", "10110010100100100100", "11000101110101001010", "00100010010011100101", "01000110010100001100", "11101101110100100111",
		 "11000010001101010101", "11010010010101010110", "00110110010100110110", "10110001010011100100", "11000110110100010101", "10100010111101100111", "11000101101101010110", "11001101111100011000", "11000101100100001001", "10110101110011101101", "00111010001100110110", "11000110011011110111", "10111110001011101010", "10111001110100000101", "11000010010100001111", "01001110111011111000", "11110110001100111010", "10110010000011110101", "00101101111100000111", "00100001100011110101", "01111110000100001001", "10101101111100000110", "00110010010100011011", "10110001010100110110"); 
		weight_ROM(5) <= (
		 "10110101100100011010", "01000110001101001001", "00110001011100011001", "01000110001100000111", "01010101111101011010", "10101101101101001010", "10111110000011100110", "00100010001100000111", "01000010110011101000", "10110010000100010111", "10111010001100101010", "11001110000100000101", "10110010010101010101", "10111101111100111000", "00111010010100111001", "11000010000100100111", "10110110010100010101", "00111010000100010110", "11000110001100010111", "01010110010011110101", "11000110001011110101", "00100101101100000110", "01111110001101001001", "00101110111100100111", "11100010010011010011", "00110010011100001000", "11001010100100110101", "11010110010100001100", "00111010000100010101", "10111010010011101000", "11000010100100001001", "11010110000011010101", "01000010001100100111", "10111110000100110101", "01011010000110011010", "10101111000011101000", "10101101000111000101", "11001010001011111010", "00111110001100000100", "01000110111101011001", "10101110010100001000", "10111110001100010110", "00100001111011001000", "00101110010100010110", "01010110011101010111", "10100101110011100101", "01001110001011100111", "11010010011101011010", "00100110100011111010", "01000110001011101000",
		 "11001010010100010111", "10111110001101001001", "11001001111101011010", "10110111001101100101", "01000110000100110111", "01000111001011110110", "00111111010011000110", "10111111010100010100", "11001001110100110110", "10111001110011001000", "10110010001110010110", "01001011001011111001", "11001110001101110101", "00110001110011101011", "11001011000100111000", "01100001111101010110", "11010001000011101000", "10100011001100110100", "00110101111100001000", "10110010010110111000", "00111010000100101000", "00101010110011100101", "01000010100101000111", "10101101111101101101", "01000110000111110100", "00110010010101000110", "10111110011011110110", "11010110010011101011", "10110110000100100101", "11001110000101010111", "10101110010100111000", "11001010100100001001", "10101010111011101001", "00111011010110101000", "10111010101100010101", "00111110111011100111", "00110111000011100110", "10111001110100101010", "10111110000110100100", "01001001100011110111", "00110001111101011010", "00111011010100010110", "01000111101011011000", "11001110001100010110", "01001110010100000101", "10101010000011010111", "10110010011100011010", "11001010001010100111", "00111010011100011001", "11000110000100110111",
		 "00101110001100100011", "01000001110101000111", "11001010000100111010", "10101010001101010111", "10111101111100001001", "11001010011100110111", "01010010100100010110", "00110110000011011001", "11010010001100010100", "01000110010011100101", "01001001111100100011", "01001010011100101001", "11100010001011101010", "10110110100100101010", "11101001110100101010", "01000101111100000111", "11010110111100101001", "10110110110101101000", "10100010000011011000", "11001010001100001010", "10111110000011100111", "00111010001011010111", "10110101110100011000", "10111110000100101001", "01001110000100010100", "01000010001101000111", "10111010001101001011", "10111101111100010101", "00100001110100100101", "10101101100100011001", "10111101110101000110", "00111010000011110111", "01000101111101111000", "10110001110100010101", "10101110001011110011", "00111010001101000111", "10100001110100011010", "00110010010100100111", "00101001101011100111", "11010010000111100101", "01001010000100000110", "01000001010100000100", "10111011001100000111", "01001010101101000101", "11010010111011110110", "00111110010100110101", "10110110000011111100", "11011010100100110110", "11000110001011110100", "00111010111011100111",
		 "11000110011100110110", "00110001111101100111", "00101110000100101001", "00110110000101000110", "01000110010011100101", "10111110001011010100", "01000010000100011000", "00100110010100100111", "01001101101100010111", "11001010010100000100", "01000110001110010101", "01000010010101010111", "01011001100011010100", "11011110010100101000", "01000010111100010111", "10101010011100011001", "01010110100011111000", "10111101010011010110", "01000010000100100100", "00111010100101000101", "11010011000101101000", "10111110001100011001", "01000010010111110101", "11010001110100000111", "11011010001011101101", "10111010011101111010", "10110110000011011001", "10110010001101110100", "01000010000100000101", "00101001111011000111", "10101010000100010110", "01010011001011110111", "10011110011100101000", "00111110011101010110", "01011010100100010111", "11001010011100010110", "11000001101100101000", "00110110010011010111", "00110001111100100110", "01000010010011110110", "11000110000011000101", "01000010001101000011", "01010101110101111010", "11010110100100111100", "01001010000011011010", "01000110011100010100", "10101110100010110110", "10110010011100111010", "11000110010100000101", "11001010001100110101",
		 "00111001111011100101", "11010010100100000111", "10111110000100101001", "01001110010011110111", "11000010011100001001", "00111010011100100110", "11010010000101101000", "00111010011100001000", "10111001111100011100", "10111010000110001001", "00100001010101101100", "10101110010100010110", "11001010011100010110", "01000110011011111000", "10111010000100101001", "01000001100011110111", "10101110010101001010", "00110001110011001100", "11001010001011100101", "00111110100011101001", "01111101110100010111", "10111001111011100111", "11000010001101010010", "00110110111011101100", "10110010011100110101", "10011010000100110101", "10101101101100001001", "00100010001101001001", "11000101110011100110", "11010010010100110111", "01000110011011000110", "01010010000101011011", "10110110010101011101", "10111110100100101001", "10111101110011110111", "00111010011100100110", "00101010000011111001", "10101010101100111001", "11000010001011010111", "00110010001101010110", "00101010111100000111", "01001011000100110110", "00100001001100100100", "01001001110100111000", "01010110000011111001", "11000010010101001000", "00111110000100100110", "10101101111100001011", "11010011011011100101", "01010010000100011000",
		 "10111010100100011001", "11000010101100011001", "10111010010100001000", "01101101110011100110", "10110110001101011000", "00111001101100001000", "01100110100100011001", "11001010001100111001", "00100101111100010101", "01001101010100011000", "11010010011100001011", "01001010010100110101", "01000010110011001100", "11000110011011100111", "10111101010100110100", "00111010010101001010", "00110110011100010100", "11100101110011110011", "10111010010100011000", "11000110100011100111", "00110110000100100110", "10111110011100110101", "11001101111100100111", "10111101100011010111", "00110110100100010100", "10100110000101011010", "00111001111100111011", "00111011010100000111", "11010010001100010101", "10110110000100100011", "01000011000111100101", "10110101111101001011", "01000110101100010101", "11001010011100111001", "10110110010100011010", "11001010001101010111", "11010010000100110111", "00110110010100001000", "01000010000100010101", "10011010011101111000", "01010111101100001011", "10110010000100101000", "11000010001100100101", "00111110100100100110", "00100010000011000110", "10101110010100100110", "01010110001011101010", "11000010001100111010", "11001010101100000111", "10111110100100111000",
		 "01000010011011100111", "01001110001100110101", "00111010111100100110", "01010101101101110111", "00110010101110001000", "00110110100100010110", "11000010111010100110", "00110010100101001001", "11001111000100000101", "10111101010100111000", "10100001110100011010", "10111101110011100111", "00110110001100001001", "10110001101100000111", "11101101110110011001", "00111010001011000100", "01100011011100100101", "00111010100011000101", "10101001101011101000", "10101001101100011000", "00111110000100001000", "00101110011100100111", "01001011000100010110", "01011001110100000100", "01000110010100100111", "11000110110100010011", "00111110011100110111", "01100010000011110101", "00101001100110010101", "01100010000100100101", "10110011000101001001", "10110010111100001010", "00101110110100101001", "01010110001100001000", "11000010000101010111", "01000111000101110110", "10110001110110000111", "11010010001101001111", "11010110101100010110", "00110001111011010110", "10110010001100101001", "00111110100100110111", "00110110110100001001", "11001110001011101001", "11011010000011110110", "10110010010101111101", "00100010001100100110", "10110110000100101000", "00101010001100110101", "00111101110100010101", 
		 "11000001111100111001", "11011110011100101011", "11001010101101101111", "00110010011100001001", "01000111000100001001", "10101110100101101000", "01000010100011110100", "11000110101100111000", "00101110010011100111", "10110110101100000111", "00111010110100001000", "01000110011101010111", "11010001111100000111", "01010110000100111000", "00110111011011011000", "11000110101100010111", "11001001110101011011", "11010010100100011000", "01010001100101001001", "01100110000101010111", "00111001101010100110", "11000110101100111000", "00111010001100000111", "00110010001100000100", "00110101110011000101", "10111010001100100110", "01001110000100010111", "00110001100111110111", "11011110000011101000", "10110110000011111011", "01001111010101110111", "00111110110011100110", "11001110010011111010", "11000010101100110111", "10110101101101010111", "11010010010100011001", "00111110010100101000", "01000011001100110101", "01011110001100000100", "00111001110100000101", "00110101101101001001", "00111110000100000111", "00101010101011000111", "11000110100101001000", "11000010000100010111", "01001010011100101011", "00110110111101100111", "00111110010011111001", "00101001110011101001", "10110010001100001011",
		 "01001010010111111000", "10110110001100101001", "00111101111011111010", "01011010111100000111", "11000101110111110110", "00110110000011110110", "01000011010100000110", "01010110011110110110", "00111001101100010111", "11001001111100000111", "01100110110100011001", "00111001110100011010", "00101001011101101000", "10110110100100000111", "11001010011110001001", "01000010011101111010", "00100001111011100111", "00111110011100001000", "10111010100100100111", "11100110001100100111", "11010110111100011000", "01000010010100100111", "11010111100101110101", "10111101110101001001", "01001110010100100111", "01101001111100101010", "01000110100100111100", "11000010000100111000", "01000010000100101000", "00110010001100011010", "10111011101100001001", "11001010111101000111", "10101101100111100111", "11011010010011101001", "01010110001100010110", "00111110000100001001", "01001001110101001010", "00111010010011000111", "11000010000100010111", "10110110101101111110", "11000010001100101000", "10110110010011111010", "11001110111100000101", "10111010001100110111", "01000010010011110111", "01000110011100001001", "11001010010100011000", "10101010101101100111", "01000001111011111000", "01010110100101110110",
		 "00111010010101100101", "01001010101110011000", "00111001101100011000", "00111010100011111001", "10110110000010100111", "01001110010100111010", "01010010010100110111", "00110010001110000111", "00101001110100011000", "00110010000011000101", "11001010000100010110", "01000001111110010110", "01001010101100010111", "00111110001100101000", "11000110110100001000", "00111001111011011000", "11010010101101001010", "10111010100100011011", "10111110000100000110", "00111101111011100111", "11000010100110001011", "11000010100100011000", "11011011101101101000", "10101110100100101000", "00111110010101001000", "11010010000110110110", "00110110101011000110", "00110001101100101010", "01000010111101111001", "00111101011100101010", "11000010100100011000", "01000101101100111010", "00110010011100111001", "01001110010011110111", "10110101111100011000", "10101010000100101000", "10110010010011100111", "00111010001011100111", "11000010100101101010", "11000010011011100110", "11011101111110001001", "01000110001101010101", "00110001110110000111", "11010110000111000110", "00110110001011011010", "01000110000100001000", "00111110111011000110", "01000010001011100111", "11010110100100110101", "01001001111100000110",
		 "00110110011011111010", "00111110000011101001", "10101001110110000111", "10110010010101001000", "10111010100101001010", "11001110101100001010", "11001010011100011000", "10110010000100000101", "10111010010100111000", "11001001110011111000", "11001010101100100111", "01001001110100001000", "00111101111011101000", "11010110101100111001", "11000101110100011010", "11001010010011101001", "11000010010100101110", "10111001110101111001", "01000010001101101001", "11001110101100011001", "01000110001100011010", "11000110100100100111", "01001010000011101010", "01000110101100011001", "01000010000110101000", "00111010011100000111", "11000110010101110111", "11010011000100111000", "11001101110100111000", "11001110101100010111", "00111011001101110110", "10111101111100010101", "10111001111100001000", "01000010011101001011", "01000010011011110110", "11011010010101011011", "00110010010110000110", "11010010011101001001", "00101001100100000111", "11001101110100101100", "01001010001100111001", "00111010000100100111", "01011101111011101010", "11000011110101000110", "10111110010100101101", "01000010011100001000", "01000011010011011000", "10111010010100001000", "01010010100100100101", "00111010000110001001",
		 "10111110000100010111", "01000010010011000110", "10111110001100111000", "00111010100011101001", "00110101111101011001", "10111010000100011000", "01011010011100110111", "01000010000101011000", "10111101111011101001", "00111110011100001000", "10110101111100001011", "11000101110011110111", "11000010000100010101", "00110010001011110111", "01011010011011100111", "01001010111011010110", "01000001111101001000", "11011110010100101000", "01000110101101000110", "01001010001011001001", "11000010010100111000", "01100010001100011010", "11000110010100110110", "10110101011100000110", "01001110001100001001", "10101111001011100111", "11000110000010101011", "01000110010011111000", "01000110101011101001", "01000110110100111101", "10110110010110001001", "11000110000100011001", "10111101110011111000", "10110110010100000111", "00110010000100010111", "00111010001100000110", "11000010000011101000", "10110010001011101001", "10110101111100010110", "11101110110100011001", "01000010010100101011", "11001010101100111000", "00101001111100000111", "00111111000101000111", "11001110010101111001", "01001110011100001000", "00111110100100100111", "10111011010100011001", "01000010001101010101", "10101001111011101000",
		 "11000010010101001000", "00111001111011001001", "01000110101101000111", "10110110000011100110", "01010110011100101100", "11000101110101101111", "00111010110011101000", "11000110011011111001", "01001011000100100111", "10111101100100001010", "00111001100011111000", "00111010001011110111", "11000010000100100111", "00111110011101010111", "01000110000100001000", "10110011000101010111", "11010110001100001010", "01010110111110010110", "10111110111100011000", "01000110110100111011", "11000110001100110110", "10111110000100010110", "01000110010011100101", "01001010000100001010", "11010010011100001000", "10111110001100101011", "11001001111100011000", "10110110011100100111", "00111001111110001001", "11000110001101100110", "11001111011100000111", "11000110001100111000", "00111110011100011000", "01000010101101001000", "10101101110100000110", "00111110011110110111", "01000010100101110111", "11000010000111000111", "01000110111101011000", "11010001110101111010", "11000001111100101001", "10110110011100101000", "11010110000101001011", "00111110001011011000", "01000010000100000111", "11001010101100110101", "11001110010100011011", "01010001110011101000", "00111110110100001000", "01100010010100001011",
		 "00111110100100100101", "01011101110100011001", "01000010010100101000", "01000101110100001000", "00110010011011010111", "01000001101011101000", "11001110000100101010", "10111110011101011100", "11000101011100001000", "10110110001100001111", "10111110011011111000", "11000110010011101001", "11011010100100110110", "10111110001100001001", "01001010001011101000", "11010010001011011000", "11001110100011010111", "00111010000100010110", "01010101111011001001", "01010110100101001001", "01010001111100000111", "00111001111100011110", "10111110001101111000", "10111010011011110110", "11000010000100110110", "00111110000011110110", "01100001111101010111", "11001101111100111001", "11000110000110001011", "01001110010011001111", "11000101111011111100", "01000010011100101001", "10111110010101111100", "00111010011101001010", "01000010110101010110", "11010101111101110110", "10111010000011000101", "01011010010100101001", "00111010010011111000", "11010110001100111000", "01000110100100111000", "01000010110100110101", "10111001010100000101", "11000110010100111000", "11011010011100110110", "01000010100101011000", "10110110000100011000", "10111101101100011000", "01000010001100000110", "11000010010101010101",
		 "01010110000100011000", "10111010011100011000", "11010011011100101001", "01001010001101011001", "01011111010101001000", "00111011001101011011", "01010110000100111001", "01000111000100011000", "01000010101101111010", "11000110100100101011", "10111101111100011000", "01000010000101011000", "11001110010101100111", "01000010000100001001", "11000010101100101001", "01000110110101011000", "11010001111100111010", "01000110001100101001", "01000110000100001010", "01000010101100011100", "11011110000111011000", "11011110010100001010", "11001110001100101011", "01100011000101001001", "11001110000100110111", "11000110111110111001", "01001010010101001001", "11001010100101111100", "11011101110101011000", "11010010010100011001", "11010011011110011001", "01010010001100001111", "01000101110100101000", "11001110111100101000", "00111110010101101000", "00111010110101111010", "01110110010100111000", "11000010001100101010", "01010010000101011001", "01000110000111111001", "11010010000100001000", "11001010100100011110", "11000110001100011001", "11010111000101001001", "01001110000101101000", "01011111000101011001", "01000110000100001000", "01000010000101011001", "01101010000100111001", "11101010100101001001",
		 "01000110100100001000", "01011010111101110111", "11000011001101101011", "01010111001101001001", "01000110111100011000", "11001010001101011001", "11001111001101011010", "01010110010100110111", "01010110011100101000", "01001011000100001010", "11011110111100111000", "01001010001011111000", "00111010010100000111", "01000110111100101010", "01001010100100001001", "11000110100100000111", "11000110100100111000", "11000010111100111010", "10111010000110011011", "01000110010100111101", "01000010001101001001", "01001110000100001001", "01001110001110101000", "00111110000101111001", "11100101110100011010", "01001010000101101001", "01000111000100101000", "01000110011100011000", "11001010010100001010", "01010110000100011001", "01001010101101011001", "10111110000100001001", "00111110001100111011", "01001110001100101000", "01000001110101100111", "01001110100100001010", "01010010011100101000", "01001110010111000110", "00111010011100101010", "01000110011100011011", "01001010001101111001", "11100110011100101000", "01001110011100100111", "01001010000011111000", "11100010110100101001", "01101010101100110111", "01001110000100010111", "01001110001100110110", "01110010010101001010", "11010111001100001000",
		 "01010010011100001001", "10111010101100011001", "01000010000100001101", "11011110100011111010", "01000010011100001000", "00111001110100111001", "10111010011101101001", "01010010110101011001", "01010110100100001001", "11010110010100011011", "10111010000101011010", "01001010000101001001", "11010011000110001010", "11000010000100101001", "01001010101100001001", "01000010011100101011", "11001010001100001010", "11000010001100011000", "01000010011100111000", "11000101110100101001", "01001010110101101011", "01000010010100001000", "01011001110100011100", "01001110100100011011", "01010010001101011010", "10111110000110001000", "01001110010100101000", "11001010000100100111", "00111111000101101000", "00111010100100011000", "01100110101100001100", "11001110010100001000", "01001110001101101010", "01000001111100011001", "01000010011101111001", "11011010111100011000", "11000110100100001010", "01001110011100111001", "01000010011101111001", "01001110001100110111", "11001010000100001010", "01001110100100101000", "01100010011100111000", "11000101110100011110", "11001110011100011000", "11011010000100000111", "11001110101111001000", "01001011111100000111", "11101110010101010111", "01000010000100001000",
		 "01001010101100101001", "11001110001101001101", "11001110010100011100", "01001110011100011001", "01010001111101101010", "11000101111011101000", "01000110010100011011", "01000110011101001011", "01011110001100101001", "01001010101100011101", "11001010010100101000", "00111001110100000111", "00111110001100000111", "11000010001100001001", "01001010010100010111", "01010110010100101000", "11000010001110111000", "01011001111101101010", "10111110001100001000", "11010001110100001001", "01001110101100101010", "11011010001101001001", "11110110101101011001", "11001010011100100111", "01010010000100011001", "11000010100100001001", "01010110101110111010", "01000110010100011100", "10111110010100011000", "00111010011100101000", "00111010001011111000", "01010110011100001001", "01010110001100111000", "10111010010100101001", "11001110011100011010", "01001010000101001001", "11010111000100111101", "11001010011100011010", "11010010011100101011", "01000110101101101001", "11101110101100111000", "01100010011100011000", "11001101111100111001", "01001010000110101010", "01001101111110111100", "01001010001100101000", "01001010100101010111", "11010101111100101000", "01010010100100101001", "00111010001101100111",
		 "01000010101100011101", "11010001111101101001", "01010010010100111010", "01000110000111101011", "11010010100100010111", "01000010101100001000", "01010010000011111011", "11000110011100111100", "01101110000011101001", "11001101111110101000", "10111010000100101001", "01000010001100111001", "01001010001100011001", "01001010101101001000", "01111010010101111000", "01001110100100100111", "11000110000100011001", "11000110100110101001", "11000010010100011001", "11000110000011111000", "11000010010110011000", "01010010010100011010", "01100110000011101010", "01000010010101010111", "01001010001100011001", "11000110001011111001", "11010010100011111010", "01001110011100111001", "11010110001100101000", "00111010001100111001", "11001110001100010111", "11001010011011111010", "11001110101101011001", "11001110110101001001", "01000001111100011000", "01001101111110001010", "11101110101101000111", "11001010000100111100", "01001101110101101001", "01000110011100010111", "01001010001101001000", "11100110010100001000", "11001010101101101111", "11001010101100101001", "11000001111011101101", "01000110001100101000", "10111110000100111010", "01000110101110011001", "11001010011110111010", "11001010110100001000",
		 "01001110000100101001", "01000010000100101001", "11001010010100001001", "01000001111110010111", "11000110010100101011", "10111110001100110111", "01010010010100001001", "01001110001100110111", "01001010010100101000", "01011010011100101010", "01000010010100111000", "01000110100110011010", "01000110110100100111", "00111010011100011001", "01001010010100000111", "01100110011100001001", "11001010010100101000", "11010011001100101000", "01001011101100101010", "10111010000101111101", "11001110000110010111", "11000110000101100111", "10111010000100000111", "11001010001101111011", "11000010011100001111", "11001010101101011100", "01001010100101101001", "11011110100100001011", "11001011000100011000", "01000010010100001000", "11000010001100101010", "01001010101100001001", "11010010001100011001", "01000010011100111001", "11010010010100001001", "11010110000101001010", "11100010001101011001", "11010010011100001011", "11000110011101101010", "11010010001100001000", "11000010010100101001", "11000110111100110111", "10111010000011111001", "01111110001100001000", "11001011101100101001", "01001110000111101000", "10111110000100101100", "11010110101100111010", "11000110001100001010", "10111010000101101101",
		 "01001010011011111000", "11100110101100011000", "01010010001100101001", "11001010001110000111", "01001110000100011000", "11010110000100001000", "01100010111100001011", "01010010001100101001", "11001010100101010111", "01000101111100101011", "10111110000100011001", "11000010000101001000", "11000101111100011000", "11001110001101010111", "11010110010101011000", "11000110110100011001", "01010110010100011001", "01111011111100001010", "11001010100100111001", "10111110000111111000", "01010110011101110111", "11001110011100011101", "01000110011100100111", "11000010011100011011"); 
		weight_ROM(6) <= (
		 "11001110000101101000", "01000110100101001001", "10111101111100100111", "01000010001100010111", "11010010001110011001", "10101110000100101000", "00111010110011110101", "01011010111100101000", "00110010011101001010", "11000101011100100111", "00110001110100000111", "01010110011011100111", "11000010010101101111", "01001110011100001000", "00111010001100110111", "01000110001100101010", "11001110101011110110", "11001010100100101000", "00110110110100010111", "01010010000011010101", "11001001111011111001", "11010101110101011000", "01001010100011100111", "00110001101100010111", "11011110000011000110", "10111111100100000111", "10111110101101110100", "00111001101011110111", "00110010001101011000", "10111110110110101100", "01000110000100110101", "00110010010011100111", "10111101110101011000", "01010010001100010111", "11001110001110110110", "10111110001100111010", "11010001101110100110", "01001110101100111000", "00111010001100100101", "00111010010011100100", "00100101111101001001", "00110011000100001001", "00111101101100000110", "10111010010100001010", "01110111001100010101", "00111010001100001000", "00110001111100001000", "00111010000011111001", "00101010010100111011", "11000110111011111001",
		 "11010110000100011010", "10111101101101011001", "00111101100101101001", "11001110101011100110", "01001001100100001000", "01000011000011110101", "00110011000011101000", "01000001111110100110", "01001010001100011000", "01000001111011101000", "10111010010100111000", "01001010100111011100", "01001001100011100111", "10101010011100111001", "11000010000011110111", "11000110010111111010", "00101001111100000110", "11001110010100001111", "00110110000101001000", "11011010101100111100", "01001110101100110111", "01000010000100000110", "11000111000110010110", "10110101110101001001", "00111001110100001000", "01001010011011100111", "11000010001011111000", "01010010010101010111", "11100110010101011000", "11011110111100111001", "01000010111100100110", "01011010001011111110", "10110101101011100111", "11000011110011000110", "01000010001100010111", "01000010000011001000", "01000110001101011001", "11001110000011000110", "11000010101100010101", "11000010111100101000", "00110001110100001001", "01010110110100000110", "10110101101011100101", "11000111101100110111", "01010010000100010111", "01000001100011000111", "01111110100100011001", "00111110100100001000", "01000011010100010110", "11001111000100010110",
		 "01000010010100000100", "00110110000100010101", "00110001100011001000", "00111110001101000110", "10101101100010111000", "11000010100110011000", "11011001101100110111", "00110110010101010111", "00111010101100110110", "00110010000011100111", "11101010010100110110", "11000010000100110111", "01001110100101011100", "10111110101011000111", "10110101111100011000", "01000010011011110110", "01100010001011000111", "10110010000011001011", "11000110000011000110", "01000001101100001000", "01100110000100001010", "01000010001100110111", "01001010001100001010", "10101010011100001000", "01001110010011010110", "01010110101100011000", "00101110011110000111", "00110010000101011001", "01000010110011110110", "00110101011011000110", "01000110110100111000", "11100110010011111010", "00110010001101110111", "00110011011100111001", "10110101110011101001", "10111010100100000111", "10101110010100100111", "00110010001100100111", "11000010011011101000", "00111010001101100111", "01000101101101000111", "01001101111100110101", "00110001110100001001", "00111010101011000111", "01000010011100001001", "11010001111011110111", "00111010101010110111", "01011101111100000101", "11001001110011010100", "11001010000011000110",
		 "01011010101011111010", "00111101110100000111", "10101001110011101000", "10101010011101011010", "01000010000100001001", "11000110000100101000", "11000010101100010111", "10111110000011100111", "00111110001100111011", "11000001110011110110", "01010010011100000111", "00111010000100001010", "01000101011011100111", "10111010001011110111", "00111110101011110111", "10101110010100011001", "10110101110101001011", "11001110011100001001", "01000110101011001000", "11001010001110011001", "01100010100100010101", "10110101111110010111", "01000010001011110110", "11001110001011101011", "01000010000100110111", "01000001101100000110", "01010111011100011000", "11000110001100010111", "00110010000011000110", "10101110110101111000", "01010010100011111000", "11001110010011111011", "11101010010100111010", "11100101101100010110", "00111010100100001001", "11000001111101011000", "11001001110101011010", "11000010100011011001", "00110010001100100111", "01101111000110010110", "00111110110011110111", "00110110101110011001", "11000010001100101001", "10101010001011100111", "11000110011100111001", "00110010010100001000", "00111010010011011000", "11000010001100000111", "01000001111011100100", "01000010001100100111",
		 "10111101100100010111", "00111010010100001000", "10111101110100001011", "01001010000011101011", "00110110001011111000", "11000010010011110110", "01000110010110111000", "00111010101101001000", "10101101111100001010", "01100110010100000111", "11000101110111001110", "01000101111011101010", "10110101110101110101", "11000110011011111000", "10111010001101101000", "11000101110011110111", "01010010001101001010", "00110010010011100111", "01000010111011101000", "11000010001100010111", "01001010000100010110", "01011110011011010111", "11010010001100010101", "00110101110100111010", "00101111011010100101", "10100110001011101000", "10110101110011101000", "10111101101101110110", "11010010000101100101", "01001110101100110110", "10111010101011101010", "10110010101100101100", "10110101110011101001", "11000001110110011101", "00111001100100000110", "00110110011100000110", "10110001111100100111", "10101101111100111011", "10111110010100011001", "00111110000100010111", "00111110111100100110", "01001010110100010111", "00101001011011100110", "00111010001011000111", "11000010100100101010", "11001101110110011000", "00101110000011100111", "10111110001101000111", "00110010001011010101", "10101010011011010110",
		 "11001011000100011011", "00110001101100101000", "11001110101100101010", "10101001101110000111", "10111001110100100111", "10110010100011101000", "00111010010110111000", "10110010110100101000", "00110110000100000111", "01000101110011000111", "00111010000011110111", "01000010011100011000", "10111010000011101000", "01010010000011111000", "11011110001110111000", "11000101111101011001", "10111010001110011000", "11000110100011110110", "10110101111100110110", "01001010100011111000", "11000110000110000111", "10110111011101010110", "11011110000100011000", "11000010110011101000", "01011110001011101011", "11000110010100001000", "11000010101100101101", "11000101101011100111", "01000010100100111001", "11011110011011100111", "00111010001101101000", "11000110011110110110", "01000010000101011000", "11000010000100011000", "10110001100101000111", "00111010001011110110", "01001110011101111010", "01101010000011100111", "11000111011100010110", "00111110010100110110", "10111110001011110111", "10101110001101011001", "11001010101100011011", "00110001111011010111", "00110010000011100111", "11100110001100010101", "10101101111100011001", "01001010000011000101", "01001010000100101000", "01000010001100100111",
		 "11001010011101000110", "01000010001100010110", "01000010100100100111", "01000110000010100111", "01001001111100110111", "00110010001101100110", "01000101100100100110", "10111110011100011000", "10111101100011000111", "10111101111010101000", "10110110000011111001", "10101010001011100111", "10111011110011110111", "01000001111100000110", "10111010011101001000", "01110110101011010101", "11000010110011111000", "00111010000100010111", "00110010011100100111", "00101001101011100101", "00111001101100000110", "00110010001100110111", "11001101110011110110", "01000010011100010110", "10111110000101110110", "00110110010011000111", "10111110000110110110", "11001010000100110111", "11001101100011100111", "01000010000100010111", "11000010010011100111", "00110111011011111000", "10110111010100110111", "00111011101100010111", "01000110010011110110", "01010101110100110111", "10111001110011000101", "01000010011100011000", "01000110011101100111", "10110110011100111010", "01010010001101001000", "00111101110100010110", "11001001010011100110", "01000001111101010110", "01000011110011110110", "01001001101100001100", "10110010001011101001", "10111110010101111000", "11010110001100100101", "00111101110100010101", 
		 "10110110001100001001", "11011010111100101111", "10110001101011001000", "11001110101011011000", "10110001111101110110", "10110010010100001001", "00111110100011110100", "00110010010100001000", "00110010000100011000", "11000001110011011001", "10110001110101000111", "11001010000100010101", "00110111011100010110", "11001110000110101001", "01001110000100100110", "11000110000100100101", "10111010001101010100", "00110010000100000100", "01000110000011010101", "00111110000011110011", "01001010111101000110", "10101001101100011011", "01011010001101010101", "10111010000011100100", "01001101110011000110", "01001110110011110101", "01000010111101110110", "11001110010100010111", "11000110001100110110", "10101011011011111000", "10111101111011111000", "01000111000011110101", "01010010010011100101", "00110001101011000111", "10110110110100010111", "10101001110011000110", "10110101000111111000", "00101110011100001000", "00110110011101000100", "00111101111100010110", "01010010011100000111", "01001110000100010110", "00101101101101000110", "00100110010011111000", "01011010100100110111", "00100110000011100100", "00100010001010100100", "01011010100011110110", "00100010010011100111", "10111110001101101001",
		 "00111110101100000101", "10101010110011110111", "01010110111011110111", "00110010101100010100", "01000010111100010010", "11101101110011000110", "10111010100011000101", "10111110111100000101", "11011010000100000111", "10111110010011101000", "00111010000101000100", "01000010011101010100", "01001110010011000100", "11000010001100111010", "01000010010100010111", "01011110110100010101", "10110001100100000110", "10101110011101010110", "10100010001011100110", "10101101110100011000", "00111101111100010111", "00111110100011110100", "10110011001100001000", "10101110011100101010", "00011011001101011000", "01001110101011110110", "11001010101100110101", "11001110000100001111", "11000001111100010011", "01110110010101110101", "10110110001110101000", "10110111001101011000", "10101111000101010111", "00111110110100000110", "00110011000100010100", "00110010011011110111", "00100110010011110110", "10110010101011110100", "10110001110100000100", "11000010010100011000", "10101001111100011000", "11001110000100100101", "00100101101011110111", "11110010001011100100", "10111010010100110110", "10100010001011000111", "00101110101100110110", "11010110001011110011", "01000011000101001000", "00111010100111000101",
		 "00110010000100000111", "00111110100101000100", "00111001101011101000", "00110110110100110101", "10110010001100001001", "10110101111011010110", "10111010100100110101", "00101101110011010100", "11000010001100010111", "10111011110011110100", "01010010001011110100", "11010001111100100111", "11000110010101000011", "10101110000011101011", "11010110011100010110", "01000010011011110101", "10111010000100100101", "10110010011011111010", "10110001111011001010", "00110010011100001001", "10110101110011101000", "01100110000101011101", "10101001110110011000", "11100110001100011000", "10101010001101001001", "10111110001011100111", "10101101101110001010", "10111101001100100101", "10110010100100111001", "10100010001010110101", "11001101110100000011", "10110110100011110101", "01000010101100111001", "10100110000100110111", "10100001101100010111", "10110001110100110100", "10111010001101001010", "10100010110100100101", "11000110101100010111", "11000111000100000111", "01010010001100000011", "00111001011100110011", "00100110100100000011", "01001001110011010011", "11000001110100101011", "00110011100101000011", "01101010000110010101", "10111110100100110110", "01001001111100010101", "10111110111100100111",
		 "01000110011011100101", "10101001100011110101", "01011110001101001000", "00100110011100010101", "00110010010011000101", "01000010001011110100", "11001110100100111011", "00101110010100110110", "10111101111100111101", "10101110100011111001", "00111001101100010100", "00110110010100000110", "10100101101100100011", "10111010100100111101", "00111010000100010100", "10100011110101101011", "10111110100100010101", "00100101010011010111", "01010110010101000111", "10100001101011110111", "01010010011100000100", "10100010000100000110", "01000110100110010101", "11011101111011000111", "01000110000110010111", "00101001101100101010", "10100101110011010111", "10111010011100100111", "00111010011011001010", "10110001100011000100", "00111110010101010100", "10111101100011010110", "10101110000100101010", "10110001111100010100", "00110110000100010100", "11000010000100110110", "01000001011100111010", "01000011011100010110", "00110101101100100100", "10111110001100010101", "00111010010011110011", "00111010000100100100", "11001101100100110111", "01000111001011000100", "10111110111011110011", "00101001110100010100", "10101110110011000100", "01000010100011110110", "01000110101100000101", "10111010010101010110",
		 "01011010000011010110", "11000101111100111001", "11000001100101000101", "01001110000011110100", "01001110110110010111", "00110110110100110110", "00111001111100010100", "00101001111101000110", "00111001111011000111", "10111101110101011000", "00101001101011100110", "11011110000111010101", "01001110011100110100", "10111010010100101000", "00111001111101001010", "10100101011101101001", "11101010000100010111", "00110011000011100110", "11100010100110010101", "11000010000100001000", "11100001110100010110", "11000010001110110100", "10111011001100010011", "00101110110110000110", "10101001101011100011", "10101010011100110110", "10100101111100001001", "00100001110100110111", "11000110011100010110", "01110110101100001010", "00101110111100001000", "00111110000011011010", "10111110111100101010", "10110110101100101010", "00101101100011000011", "01000110011011110101", "00101010101100100111", "00110001110100111100", "11001101110100010110", "01010110000100001000", "00101010001101000111", "10111111001100110111", "10101001011011000011", "11001110011100101010", "01000010001100001010", "01001010101100110101", "11000001110011110111", "10110110011100111011", "11001110001011110100", "00100010001100110110",
		 "10110110001011101001", "10111001010100011000", "10111010000110001000", "00100010001101000111", "00110101001011110101", "01000010000110001001", "11001110011110000111", "11000101111100011001", "00101101100011100101", "00100101000010001001", "00111110100011110111", "10100110100100010111", "10110010010100101000", "11000010000100100110", "10100101010100010101", "10110101110011111000", "00111010011100010110", "10111010000110110110", "10101110111011000110", "10110010001100010011", "00101010100110000110", "00100010111100010100", "01000001101011000101", "00101010001100110110", "11000010001100100011", "00111110110011111001", "10110110011011110111", "10110101111101100101", "01001010010100000011", "11000110011011101011", "11001010111100110101", "11001010011100101001", "10111010011100100101", "10110110000100011000", "10011011010100000111", "00111010001100001000", "01000010000100011001", "10101110011011100101", "00111110011100010101", "10101001100011100100", "11000110010011111010", "00101010011011001100", "00101001010100100101", "10110110111101000110", "00101010010100000110", "00100110001100010101", "01010110101100011000", "10111110010011000011", "01000010011100000111", "11001010000011110110",
		 "01001010001011000110", "10111010001100000011", "00110001111100000111", "10111101110011110110", "01001010101101010101", "10101101110011100111", "11001001110101010101", "00110010011100000101", "00100101101100000100", "10110101011100101101", "10110110011011101100", "10110010001011101000", "10111010011100001110", "00110110001101101010", "11000101101110001101", "00011110101100000011", "11000011111101010101", "00101110010011100101", "00110001100100100101", "01001001100100000111", "01001110010100110110", "00110010001011000110", "10110010010101010110", "10111001110101001000", "10111101110100010100", "00111010001100110011", "00101010000100010110", "01000001110011110101", "01000001001100110101", "00101110000101100111", "10111101111010100110", "01001110010100001010", "10101110001100100110", "01000010001101001010", "01000010000100111001", "11000101101110110100", "10111101111100101010", "11010110011100011101", "10110110100100010011", "00111001111100000101", "11001001111011100101", "00111010000101010010", "10111001100100000110", "00111110010100110111", "00111011110011010110", "10101001111100110100", "00101011101011110101", "10111010010100001000", "00110001111100100110", "00110010100101011001", 
		 "10110010011100001010", "10110101111011000111", "10110110011100011001", "00111001111100100111", "10101011101100111000", "10100110001100000111", "01000001100011110100", "10110110100011111001", "00101001110011000101", "00111111011100100110", "01010001100100000110", "01011101110100110101", "01000001110011010111", "01001001111011101000", "00110010001011110101", "01001101111100010101", "10111010001101010011", "00111001100011010111", "00110010010100110110", "00110111100011010110", "01111001101010111000", "10111110110100010111", "11010001110100110111", "00110001101011001001", "01000101100011100100", "10110010000011000100", "10111110001101110100", "00110001110111110101", "01000010000011010110", "10101110100011101000", "01001010011100010110", "00111001110011100110", "11000101101100010110", "11000010000101010101", "10111010111100011000", "10111110010101011010", "00110101100011111000", "01010010001100000111", "00101010001011100100", "00101010000011100101", "00110001101011000110", "00111110010110001001", "00111101111011000110", "00111010001011100111", "01010010101100010110", "11010001111101111001", "00100010101011100101", "01000001100011010110", "00111001100011001000", "10101110001100000110",
		 "01111110011011110111", "10101101111100001000", "00110101101011100100", "11101010001011100110", "11000001011100011011", "01000010100010110101", "00111010010100011000", "10111110001101110100", "00110001101010100101", "10110001011011000111", "00110010010110010101", "11010010101101010110", "00101001100100000110", "10101110110100011000", "00110010101011110110", "11000110010101110110", "00100001000011000100", "00111001110011100111", "01000110010100011001", "01000101101011111100", "00111010100100110111", "00101101110101010101", "01010101110011110110", "10110110001101000110", "01001001010010110110", "00111010101100011001", "11000001111011110111", "10111110010110110111", "10111001110011110110", "01000001111011010111", "00111001111100000110", "10111110000011010111", "10101101111010101001", "10110010011101110111", "11001001101100000110", "00111001111011011000", "01000010000011000110", "01000111010011110110", "11000001111100011010", "10110010101011111001", "11001110110011110111", "00111001101100000111", "10111101111100000101", "01000111001101010110", "01001010000100010110", "00101001011010100101", "10100001110011000111", "10110001100100010111", "01000010111100110110", "01011001110011110101",
		 "00111001111100000100", "00110110000011100111", "11001001100100100110", "10111001110011100110", "10101010000010101000", "10110110001101110110", "11001001111100110101", "00100001110011001000", "00110001111100101001", "00101010000100000100", "01000010011011110100", "01011010000100010110", "00110010101011100111", "00111001111100001001", "10110101110101110111", "00111010001011010110", "00111001011011011000", "10110010000100101000", "10110110011100000111", "00111001111011001000", "00111110001011011001", "00101010001100100111", "11001101111100000111", "11000111001100001000", "00111001110100100101", "01001010011011110100", "00101101101110000111", "00101110001011011000", "00110011110100010101", "01011001111011000111", "01000010010100001111", "00110010000011010111", "00101010011100010111", "11011001110100010100", "10101101010011010110", "10101001010011111011", "10110101101011101111", "10111001101010101010", "10111010011100011001", "00111010000101000110", "10111001110100100101", "00110001111011110101", "00101001011110100100", "00100001101100000110", "01000111101011110111", "00111010001011010111", "01000011111011110101", "01111110001111000100", "01000110100011010100", "10110110010011000101",
		 "01001001111100111001", "00110010010100000111", "10101001010011100101", "10100001101011000110", "11000101100100010101", "11000101111100110111", "11001110000100110110", "11010010000100001000", "01000110001100110101", "00110001100011010101", "00110001101010100111", "00111001100011000111", "11011101111100000110", "10111110010100101011", "00110110001011100100", "10110110100100011001", "10101110000111111011", "01000101100101101110", "00100001111011000101", "01011110011100011000", "00110010000011010100", "10110110000011010110", "00110001111100110110", "10110101111011011000", "10111011000100010111", "10110010011011000101", "01000101010011111000", "01000110001100010100", "00110001110011101001", "10100010000010100110", "01010010001110110100", "10101101010011100111", "10101110010101001001", "01000101101010110101", "00110010000101110101", "10110010001100001000", "00110001100101000111", "10111001110011111011", "00110001110100111100", "10110101100100110101", "00111001101011011001", "00111011000011100111", "10111110010100101000", "10100010111100100100", "01000010010011011000", "10110001111011111000", "00110001100010110100", "10101101110100101000", "00111101110011000101", "00111110001100010110",
		 "11000110100101110101", "01000010000100110100", "10101110001100011001", "00110010001100000101", "00111101010011101001", "00111010000101000111", "00111001111100110101", "00101110110101011011", "10101010000101101011", "10110010011110100111", "10110101110110101000", "00110101101011000100", "10111010011100110101", "11000110011011001000", "10110010001100000110", "01000010010011010110", "10111001010011001000", "01000010000011110110", "01111110011011111001", "10111010101011110101", "10111010100100110110", "11000010111011001001", "10111010000011010100", "10101101100011101000", "00110010001011000110", "10010001100100011010", "10110101100011100111", "01001101011101010100", "11000010010100010111", "10110101101100110100", "00111010000100000111", "11000010000100010111", "10101101010011011000", "10101110010100111001", "00101001110011000101", "00110001100011100110", "10110010011100001000", "10100110001100000110", "11000101100100010110", "00110010000011010110", "11100001101011000101", "11001001110011110101", "11000110001011000101", "01000010101011001000", "10111101101100110111", "01001110100110101000", "00110101110011000111", "10110101110100011000", "00100001101011110110", "10110010011011001101",
		 "10111101111100010111", "10101101011100001000", "01010110001100000111", "00101001011011100101", "00100101110011000101", "01011110011100010111", "01000010000100011001", "10111110000101011000", "01010110011100000111", "01010101010010100111", "00110010000011111010", "01100010100110110101", "11000001111101100110", "10101010001101101001", "10110101100111010101", "01000001100100000111", "10101010011100110100", "10100101010100010101", "10110101110100110110", "01001001110011110100", "01000001110100010110", "10101110110100010110", "00110101111011110111", "01001010000010111101", "10111011011100010110", "10101010011011100101", "10101101111100101010", "01001010011011100111", "00110001111100000011", "11001010111011010101", "01001010101011110101", "10111010100100010101", "01011110100101000111", "10110110000101110111", "10111010000011000101", "01001110000100110111", "01000101110100110101", "00101001000011000111", "11011110001011110101", "01011010010100010111", "10101101111011110111", "10110110111011000111", "11011110010101100110", "01000010111010110111", "00101010010011000100", "10110010101011011000", "10110110101011001001", "11000001100011000100", "01001010001100101000", "10101001110100001000",
		 "10110110001011000110", "00110110000101010011", "01000010101011110110", "00101101010011000101", "11001001101011100110", "00110001101011000110", "00111001110010100111", "10111110100100001001", "00110101000100100100", "10101101101011111011", "10101101110100010111", "10110010100010100111", "11001101111011000110", "00110001101011100110", "10110110001100001000", "00111010101011010101", "11001101101100110111", "10111111010011011011", "01001101100110000110", "00011001010011100110", "01001001100101011000", "11001001111010100100", "01000101010011110111", "10110110111011110101");
		weight_ROM(7) <= (
		 "11000001110101011000", "00111001101100000110", "00101001010011001001", "00111001111100000111", "11001011110100100111", "01000110001011101000", "00111001110100100110", "00101101110100000111", "10110110000011001001", "11001001110100101101", "10100110111100011000", "11001010100100111001", "11000010001100000110", "00110010101101010110", "11010010110100111000", "01010010000100101000", "10101110101011100111", "10101010000100000100", "11010110000100000101", "01000011010101010011", "11000010011100010110", "00100010011100100101", "01000110011100111010", "10111001111100100101", "11001001100011110100", "10111110101110010101", "11010010010101110111", "01000011001100111010", "00111101111100010100", "01010010111100111001", "11010010001101000110", "01000110100011000101", "00110010000100001000", "11010110111100000110", "10111110100100111001", "00100101100011101010", "00101101111100101000", "01010110001101100111", "10110001111100100011", "01000010000011100111", "00011001110100101001", "01000110001100010111", "10110101101101000110", "10111010010011101000", "01010010000100011000", "00111110000100000101", "01000110010011111001", "01010101110100000110", "00101010000100010111", "10111010010100101000",
		 "11100011010011110111", "01001001011011101001", "00110001011100000100", "11000001111100100100", "01001111000100110111", "10110010000100000101", "11000011010100110100", "10111001111101000101", "10100110001101101011", "11001011000011111001", "00110010100111010110", "11000110000111011000", "01001001011101010101", "10110010101100101011", "01000010100011110110", "01000010100111010111", "10010110001100001000", "00110010001101110011", "11000101011100111000", "10110110001011011000", "00110010000101011000", "00101010010011000100", "01000010000100101001", "01001010010101001010", "11010011110101010111", "01001010010100110110", "01001010000100110110", "01000110010100111010", "01001001110011100111", "01001001111100010111", "00110101110100001000", "11000011111101001000", "00101101111011101100", "11010010001100110101", "00111110011011100100", "00111001100011111010", "10110010110100000110", "01000010001100000101", "11000010110100110101", "01010110000100111000", "10110001010011111000", "00111110100100011010", "11000010100100110101", "11010110001100110110", "11000010011111010111", "11000001110011000110", "00110010110100000110", "01001110010011100011", "01000110011101011000", "00111010000011100100",
		 "00110010101011110111", "01111101110101011000", "11000010111100100111", "11000011001101110101", "10111001110010111011", "10111010111011110110", "00111001111101101000", "11000010011100011000", "11010010000011110101", "00111010000011000101", "00111111000100010101", "00111010011100011010", "11001110111100110111", "10111111101011111010", "00111110000100111000", "01001110000111010111", "11000010001011001101", "11011010011100111001", "10100010000101001000", "10101110000100101010", "10111110000011010110", "10111110010101010100", "10110110100100010111", "10111010001100011000", "01000111001100010011", "00111010000100100100", "10110010011100101001", "11011001110101000111", "00100010010101000111", "00110101011100111001", "10111010000100010101", "11100010000011110101", "01100110001100111010", "00110010010011110101", "00101101010011000101", "10101110010101000110", "10100101011101001000", "00101010001011110110", "10111001110100000111", "00110110000100110111", "11000010001100010101", "00101001101100000100", "10111010011011100110", "11001011000100101000", "01011110110100110101", "10101010010110100101", "00110001101011000100", "11110010000101110100", "10110010010011110110", "00101101101100110101",
		 "00111110000100101000", "10101101101100101001", "11000010010101101001", "10100010000100110101", "10111010010011100101", "10111110101011110110", "01000010011100011001", "00110010000100100110", "01010010000101011000", "10110001110100000110", "00110110001100000110", "10111010011100000110", "00101101111101100100", "11000010001011100111", "00110010101011110101", "10111010010100011100", "11000010111100011001", "10111110000011110111", "01000110011101010111", "01000110011100011010", "11000110011101110101", "10101110010100001010", "11000110110100110111", "11001110111011100110", "10110110000111110111", "10101101111101111001", "00100001100010100111", "10111010010100010111", "00100110010010110111", "01000001101101000111", "11001010001110010100", "01001101110011101001", "00111001111101000111", "01000001111011110100", "10111010000100110110", "10111110101101000110", "01001110101110111000", "01010010110011100100", "10110010001101010101", "01001001111100110101", "00111010110100010110", "01000010011011100110", "10110101101011110110", "11100010110100011010", "11011110010011110101", "10110001111100101000", "10111110010010100100", "10101001110100101000", "00111110100011000110", "10110010001011010101",
		 "01001110000100111000", "01001010100100000100", "01001001111100111100", "01001010010101100110", "01010011111101110101", "10101001110100100110", "01010010001100011000", "00110110011100001000", "10110110100011100111", "01000001101100111000", "10111001101100101000", "00111101111100000110", "01010110001100110110", "11000110011011101000", "10110110001100100111", "11001001110101010101", "10110001110100100111", "11001110010110110110", "11011010010100110110", "01010010000110101001", "10111110011100010111", "01100110101100111000", "00111110100100110011", "10100001100100101000", "01001010011101110111", "10100101111100010101", "11100001111100011001", "00111001100111010111", "11000110001101001001", "01001010011100010111", "10110110010011010111", "01100110000101111010", "10111110001100101001", "11100001111101101001", "00110010010100110111", "10110010101100100110", "00111010000011001001", "10110110010100111000", "10111010100100111101", "11101010000100100111", "00111001110100100100", "01000010001100010101", "00110101111100000111", "10111010001011010101", "11000011001100110111", "00111010000100000101", "11001101110100010110", "10111110010110111011", "00111010001100000101", "01000110000100111000",
		 "01101011000100111011", "00111101100101000111", "11001101011101001000", "11000110000100100110", "00101001101100101000", "00110001101100100111", "10111101110100001010", "00111011011011100111", "00100101110101010101", "11000101110010110110", "10111010101100011001", "10111010011011011011", "00101101110101101000", "11010010010100001000", "10101101110100010101", "00101111100011111011", "10110110001011111000", "10110110001101000101", "01001010010111111010", "00110010000101010101", "00111010111101010111", "10101110100101001011", "00110101110011010111", "01010110010011010101", "11001110010101010110", "11001010000100001001", "00101001110100001000", "00101001100100110110", "11001010010101010100", "01000110011011100100", "10111110011100010111", "01000010001100110100", "11010001111011110101", "01001111000100100111", "00101010000011000110", "00111010101011110110", "01001010010011110111", "01000001110011110101", "01111110100100010110", "10110010000101000100", "10111101111100010111", "10110010011101011011", "00110010110100101001", "01001010010111010110", "00111110010101100110", "01000110000101100101", "10110010010100001001", "00110111001011100110", "01001111011100101010", "00011001111110011000",
		 "00111101110100010101", "01000010010110011000", "10101110000100110111", "10110101010100010100", "11001010001100111010", "10110110101011101000", "11001111010011110110", "00110010011100101000", "01100101101100101000", "00111001111011101010", "10100110011100100111", "10111010110111101111", "01001010011101010111", "10101010100101100110", "11010110111100110111", "10101110001011100101", "00101001110100100110", "10101010001100000101", "10111110011100101000", "10101010111011101000", "11001011010100101000", "00101110011100000101", "00100001110011111001", "11000001101100000101", "11000010100011110110", "01000001111100010100", "10111010001100001000", "10111110100100000110", "00101101010101010011", "11010110010100111000", "10110001100100100111", "00111010011110010111", "00101010100100000101", "11000101110011111001", "01000110010101110110", "01000110000011110110", "10110001110100010100", "11001010001100011000", "01001011000100100110", "00110010101010110110", "00110010001100100101", "11101010011011100110", "10111110110011100111", "00110010010101010111", "01001110100100000110", "10111010000100011000", "11001001110011100101", "01010110000100010111", "10110110010100111001", "00111101110100010101", 
		 "11010111000101000111", "01111001101100111001", "00101001011011110111", "11001010101011100110", "01000010110011100110", "01000101110100101000", "00110110010100010011", "00011110000011101000", "00110101110011100110", "10101110100100110111", "00110010001101100111", "01000110100100100100", "00101001101011000100", "01000010010101010111", "00111011001100100110", "11001010110100010110", "01010110101100110101", "01000010011100001001", "10101101110011110100", "11001010100100010100", "01010101111100100111", "10100101111100101000", "11010101110101000111", "00110111001100100100", "00111001010011010101", "11101110010011110101", "01000011010011110101", "11000010010100010111", "10110010101100010111", "10111010011100000111", "01001010010011100110", "00110110110011100100", "00111010000110000100", "00110010001100010111", "10111110011100110111", "10110010010011000111", "00101001110011111011", "01000010011100100110", "10110001110100000101", "11000111100101010110", "10111001101101001000", "01000101111101110100", "00110101110101001010", "00101110000011010111", "11010110001011110111", "10101010101011111001", "10111110011100000011", "01011001110101110111", "00110010010101101000", "10110010011100101011",
		 "01000010010100011011", "10111010011101011010", "11010001101100010011", "00011010011011100101", "00110001111100110101", "00110010001100000100", "01001011010011101000", "10100110001011100100", "01000110101100111100", "01100011000011100110", "00110010010101000011", "11001010000100110110", "01000001100011100110", "01000010010100000111", "01000110010100110110", "10111010000100110110", "10101001100100101001", "10110010000100110100", "10101101101011100110", "10110010010100101010", "11100010000100110101", "10110010001100110110", "10110101110100101000", "00111110000110000111", "00110110011101010101", "01010011000100111000", "11000010000100010101", "11011110010100010111", "11000110101100010100", "11011010010111110110", "11000101110100101100", "11001110001100101000", "11001010111100110101", "01001111011101110110", "10111111000100010100", "00111110100011001000", "00110110101100110101", "10101010101100010101", "11010101110100010100", "11001110110101111010", "10011001100011111000", "11001010101100100100", "00111110001011010111", "11011010010011110110", "00110101110100011001", "10100110001100010110", "00011001110011000111", "10111101110011001000", "10111010001100111001", "01000010000101000011",
		 "00110101110101001000", "01000001111100110100", "10111001110100101000", "01001110100011110101", "11001010001011000111", "10110110000011110111", "00110110010100011001", "00101010010011100111", "01010110000101111001", "00101010000011110100", "11010010001100001000", "01001110100100110111", "11011010001100100110", "11001101110011011001", "10111010010110001001", "01000010110100110101", "01001110101101010111", "01011010011100001001", "00101110010101001001", "00101110101011101000", "10111110001100110111", "01000110011101110101", "10100010011011110110", "01011010011100100111", "11000010100011100110", "10111010010011100100", "01010101010100100111", "11001101111100010101", "10110110111100100100", "00100101101100010101", "01000010110101000110", "00111001110011100100", "01000110010101011001", "10100010000011100101", "10111101101100100110", "01010010011100010111", "00111110101100011001", "10110110001100110111", "11010010010100011000", "01000010011100000110", "01101001011100000101", "00110110111100010110", "10111001111101100011", "01001110000100010110", "11000010011100100101", "00110110011100111000", "00110010010011010101", "11000110011100111001", "11000010001011110101", "10110110101011111001",
		 "01000110101011010110", "00111010000011011100", "00110110110100100111", "10101110000100110110", "00111110000011100100", "00110101111010100100", "00111110110100010110", "10101011010011001000", "11000110010100110110", "10101010000110100101", "00111101101100010110", "00101110000100101000", "10101110001100100100", "10110010100100101010", "01001010010100010011", "10110011000101001001", "00111110110011101010", "10111101101011110111", "10101001110100000110", "10100110000011101000", "01111001110100010110", "00111010001011011001", "00110111011101110101", "11011110010100111001", "01001010101100001110", "10111111000101001010", "00110001010011101010", "10101110011100100110", "10110001111011100101", "00110001100011010100", "01001010101100000101", "11000110001100110110", "10100010000100101010", "01010010001100010100", "10111110010011100101", "10110010011011110101", "01001001100011110111", "10111010001100110111", "10110101100011000101", "01010110000100110101", "00110110010010110100", "01001010100101111100", "10111011000100111001", "11010110001011000110", "11100010001010010110", "10110011111100010101", "00110110010010000011", "00111001111100010110", "01000110111100000110", "00111110010100010101",
		 "11000001111100001010", "00110010010011000100", "10100001101101011100", "01010110001100010101", "10111110110011110100", "11010001111100000101", "01001010000011110110", "00110111000100000111", "00101010001010100111", "11001010001100001010", "00011001010100111000", "11001110000011010011", "11001010100101110101", "01000111000101101001", "10100110110011011001", "11001011011100100100", "00110011010100000110", "00110110111100010100", "01000010111100010100", "00111001100011111010", "11000110000011111000", "11000110110100110110", "11011010010100010011", "10100110000101100111", "10100001111011010101", "10101110010100010101", "10011101111100000111", "01000001011011010100", "11010110000100110111", "10111110011011101000", "10110110011011000110", "01001010011100001000", "11000010011110011000", "10111010000100111010", "10110101100101100100", "01000010111011110101", "10110111011011111001", "00110001100100111001", "10110101111100101001", "01010101111101100101", "00111001111100100100", "10111010101111011000", "10011000110100000110", "11000011000100011010", "10110110010101001011", "11000110010011110110", "11000001110011010011", "10101111000101100110", "11011001111100110011", "00110110000100110110",
		 "11000110001011110111", "00100101111101000111", "01000110011100001000", "01010001110101001010", "00100101100101011000", "11100011010100100110", "00111110011100000111", "11011110101011111011", "11010001010110000100", "00100101101101011001", "01100010101100011010", "10110010101100000101", "10101101110101001000", "10111010010011110110", "10101101010100000110", "00111110001100011001", "11001110100100110100", "01000010101100000100", "10110010011100001010", "10110010011101100111", "00111010110100000111", "00101010011100000110", "00100110000011100110", "00110001000100111010", "11001110101011000101", "10110111001111000111", "00111010001100101001", "10110101011100000111", "11010001111101100101", "10101010101011100010", "11000010001100110101", "10111110100100100100", "01000110110011100101", "11010110001100000111", "10111010110101010111", "11010010100100111010", "11001010011101111011", "00110111001101000101", "00110010000100110110", "00101001101100000101", "11001011101100011001", "00101110101110110111", "10111010010101011010", "00110111101100100100", "10110111001100100111", "10110110001100110011", "01100110111110010111", "00111010010011000111", "11001001110100001001", "11000001111100000011",
		 "01000101111011110110", "01001010011100000100", "00110110111100010110", "11000001110100011000", "01000010001101010100", "10101110100100001000", "11000110001011011000", "00101010101011100110", "00110110001011100111", "10110101100100101010", "10110001111100001100", "10111101111100011000", "10111010000100011010", "01011010000100000111", "10111110010101101001", "01000010001011010110", "01000110110100000011", "10111110110011000110", "00110101011100000111", "10101001010100011010", "01000011100101001001", "01000110101011000101", "10101101111100110101", "11000010101011100111", "10111010001100110100", "00110110001101010101", "00110010001011101010", "11011001110100100100", "00100001010100010101", "00111001110100010101", "10100110001100111010", "11000010001100111000", "11000010011011101000", "01000010101110000110", "00111010101100110101", "01000010010100110101", "10101010011100011000", "01010110101011111001", "11010110000111001000", "10110010011011001000", "00110010000010110100", "00111001110100110100", "01011001100011110110", "11001010001011111001", "01000110100010100101", "10101110010011110101", "00111110100100000100", "10110110101100001010", "01000010010100010100", "00100001101011000101", 
		 "11010110111101111010", "10110110000101101001", "01001110000011111001", "00110001101100000111", "01001010101100001001", "10101011001100000110", "00111001110101010101", "11001111000011101000", "00101010000100000110", "10111110010100110111", "00111001100100001000", "01010110110110110101", "10111110101100010111", "00111010011100100111", "00111010001011011000", "01000010010011110111", "11010110001011110101", "11000110110100000111", "00110010011110010110", "11010110101100010101", "00110001111010101000", "11100101111011011011", "11001110011100100110", "00111010001011111001", "00111010110011101000", "10110010000011100111", "10111110001101110100", "00101001110100010111", "11011011110011011000", "10101110010011001001", "10111110001100010101", "00110010110100111010", "11001101111100110111", "10111001110011110110", "11000101111011110111", "10111101110011110111", "01000101111100100110", "00111001110111011001", "01001110101011000110", "01010010000011000110", "00101001101011000110", "00111110100100001001", "00110101101011101000", "10111001111100100111", "11001110000110011000", "01001010001100111000", "00101001101110100101", "01000111100100110110", "00101001110100001000", "10111110001100001001",
		 "01001110010101010110", "10111010011101011001", "01001101111100000110", "10111010111100000111", "10111001111011110111", "01000101110100010111", "00111010010100000111", "11000010011100010110", "10111001111010110110", "00111001111100001010", "11100011000100110111", "00111010001101011100", "00111001100100000111", "10101101110101011001", "01001010010100010101", "01100010001100101000", "00101001001101000111", "01001010000101100111", "11010110010101101000", "01001101110011111000", "01011010010100111001", "00110010110100101011", "11010101110011110110", "10110101100100101000", "01010110110100001011", "00111010001011101000", "11001110010011011000", "11000110011100011000", "01001101111101011000", "01000110111100011000", "00111011111100101000", "10111110001100101000", "10110101111100000111", "00111010000011101100", "01001101111100111000", "00111110001100101000", "01000001110100100101", "01101010110100011001", "10111110110110010111", "10111110010101011001", "10111010101100011000", "11000110010100100110", "11000101101100000110", "11001110100101001001", "01011010001110101011", "00111110110011000111", "10101011111100011010", "10111010100011110111", "00111110101011010111", "11000110010100110101",
		 "00101001111100100101", "00101110000011011000", "10110001100101101010", "01001010101100111100", "10110001110011000111", "11011001111100010110", "11001010001100110111", "00100010000011100100", "01000001110100101001", "00110011000100000111", "00111110000011110110", "01010110111100110111", "01000001110100011000", "01000010111111000111", "10111110011101011001", "01000001101100110101", "11010001101011101000", "10100110000010101000", "01001010000011101000", "00101110011011001000", "10111001110100001000", "00110110001100101000", "10110010100100011100", "10111110110100000110", "00111110010100000101", "11000010001011010101", "00111110011101100111", "00110110000100000101", "00111101110100110110", "00111101011101000110", "01000010001100111000", "01101101110100001000", "00110001111100001111", "01011101110100010110", "10111110000101010111", "10110110100011100110", "10101101110011111010", "00111010101011000110", "10110010000011111011", "00111001110110000100", "01001101110100100100", "01100110001100010101", "00101010000100000110", "10110001101100000110", "00111110001011101000", "00110001111100000101", "00110110011011110110", "11100101111100000101", "01001111000011110110", "00111010001100000101",
		 "01011101111100010111", "00110110000011100111", "10111010000110100111", "10100011011011100111", "11001010111100010111", "10111110001011100101", "00111010001100110111", "11001010000100101000", "10111010111100010111", "01000010010011110111", "00111010010110011010", "01010001100100000111", "00111101101011001000", "10111010011100101000", "01001101110100000101", "10110010100101011011", "10111110011101001000", "11000010111100000111", "00110101111100000110", "11001110101011111000", "01010010011101010110", "01010011110101010111", "00111010001011100101", "11100101111100111010", "10101101110011101000", "00111101111011100111", "10110101111011111000", "01100110010100110110", "11010110011100010101", "10101010011100010111", "01000010001100010110", "11000101100011011010", "10101010001101011011", "01000010001100100110", "00110001100100010110", "01000001101011101000", "01000010000100000101", "10111001100100101111", "00101011001110110110", "11010010011100101010", "01000111100100000110", "00110010000011010101", "01100110001100101000", "10110101110100110110", "01100110101100100110", "10111010100101000110", "00111001110011110111", "11001110001101001000", "01010010100011100100", "01000010001100100110",
		 "10111010111011110101", "01001111000100000110", "10111110100011111001", "01000010000100100111", "00101110000100010111", "01000001110101010101", "11011010011100110111", "11001010001101111001", "10110010000100001010", "01111110011101100111", "00110010010101001010", "10111110001101101011", "10111110000101010101", "00111010001011001011", "10101010001110101010", "11011010101100110110", "00111001110100001000", "01000010010011000110", "11001110010101110111", "01001010001011111000", "01011010000100001010", "11010010001100100110", "00111010010100010101", "10110101101100111001", "00111010101011000110", "10100110100100100111", "11000110000011100111", "01111010011100110111", "11010010101101011000", "11001011000100111010", "00111001110100101001", "11000010011110001001", "10101101110100010111", "10111110010011101010", "00111110001101100110", "01000001111100000101", "10110110101100000110", "10110101100100101001", "10101101100101010110", "00111110000011101100", "10110111011101000100", "11100110011100110111", "11001101011011100111", "00111110011011100111", "10111110000100001001", "10111010011100110101", "00111110000011100101", "10111110100100001001", "00111010000100000111", "10110010001011110111",
		 "11001010001100101010", "10111101111011100111", "01000110011101100111", "00111010001100000111", "00110001101101100110", "11010110011100101010", "11101010000111101111", "10110011001011111010", "01111111000011000110", "11000101010011011100", "01000010010011001010", "00111010010100110101", "10110110000101001000", "10110010011100100111", "01100001111101111001", "10111101111100111000", "10111101111011110110", "11001101101101110110", "10110110000100011010", "01000111000100100111", "01001110000100010110", "10111010111100110111", "00111010010011110111", "00110010110011000111", "01011110011100111001", "10110110000100001011", "10111110010100101000", "01100110101011000110", "00111110011101110111", "11000010011011101001", "00111010011100110110", "10111101110100010110", "01001110010101110110", "11001001111011110111", "10110110010100000100", "01000010011100011000", "01000010010110011010", "10111001100011101001", "11001001111011110100", "11010010000011110110", "11000001111011111000", "10101010001101011011", "11010101110011111100", "00110010011011011001", "00101111000011100110", "11001010010100010111", "11001110000100111001", "11010001110011100110", "01000010011100000111", "11000010001101000110",
		 "01000010111011100101", "10111010101101110101", "10111110010101000111", "01000101100011100100", "01011010011110010110", "00111010101011101000", "01010001100011000110", "10111101110100001000", "11000101000011100110", "10110110001100111010", "10101010001100111010", "10111101110010101011", "11010010000100010110", "00110010001100000111", "11001001111011101000", "01001101111100010111", "10111010101110110111", "01001010010011111010", "11011110000101100110", "00110101111100000110", "01001001100100100111", "00111001111100100111", "01010101100011001001", "00111001101100010110"); 
		weight_ROM(8) <= (
		 "11001110010101111000", "01011010110100011011", "11001010001011101000", "01001110011100011000", "11010110101100000111", "10101110010011110111", "11010010000011101000", "00111010000100001011", "00101101110011111011", "11010001110100001000", "10110110010100011000", "11010110110111001000", "00111010011100000100", "01001010010011111010", "01001010001101111000", "01010010110101001000", "11001010011100111000", "01000101110101011010", "11000110010100000101", "11001110000100010101", "10111010100011110111", "01001010011100001001", "01001110110100001001", "11000010000100111011", "01000010011100010110", "00111111100110010100", "01000110000101001000", "10110010010100101001", "01000010101011010110", "11000110010100011000", "11011110100011111011", "01000010000011100101", "01010110011011100101", "11001110010100001110", "11001110010100101001", "01000010001100011100", "00111010010100101000", "01100110101101000101", "11011110010011100111", "11000110011100100111", "01011110001110101010", "11000001111101101000", "11001010001101011000", "01000110111100010111", "01110010010100111000", "11000011001100000110", "01000010110100000111", "01000010111101101001", "00101110001101011000", "11000101110100101001",
		 "10111110010101001010", "01011010110011101010", "01101001111100110111", "01000110011011100110", "01000110110101111000", "01000101110100010111", "11000010000011101011", "11010010010100111000", "11000110101100101111", "11001010010100001011", "00111010000100101011", "01010010010100101000", "10110110110100110110", "10111110100111111010", "11010010010101011010", "01010101110100010111", "10110101111100001001", "01001010010100010100", "10111011000100101001", "11000010001100111000", "01000010010101001010", "11001011111100100101", "11010010111100111001", "01000111000100000111", "01010010011100110101", "01000010011011101011", "01000110001100110111", "01000110010101011010", "01010110100100011001", "01000010000101111101", "11000010101101101000", "01010001111011101001", "11000110001101101000", "11010011010011101011", "01011110110101000110", "11000010010101111011", "11001011010100000101", "01100001111110001001", "01001010010011111010", "11010110010100000111", "01010110101011001000", "01010110011101100101", "11010010111100000110", "11000110011100010110", "11100110101011101001", "10110110000100011011", "00110110001100011001", "11001010010101000111", "00111110110100111000", "01000001110100100101",
		 "01001010011100110101", "10111010000101101000", "01010110011101001001", "01000010101101010111", "10111110000101111000", "10111110001100001100", "00111010000101111000", "11001110100100000111", "01000010011100010111", "11000010001100100100", "01000001110100100110", "01000010011100101011", "01010010000101000111", "10111001110101011001", "11101010011100000111", "01001110010100000111", "11001011001100101111", "11000010000100101000", "10110110110100001011", "01000110100100001000", "01001010010100101001", "11000110010100110110", "11011110011100001000", "10110110010100110111", "10111010100100100111", "11000110011100100101", "01000110010100111001", "10110011001101000110", "11000001111100001000", "10111110011011100111", "11010110001100111000", "11000110101110110111", "01101110101100001001", "11011010000100000101", "00111001110011111000", "10111101110101001000", "10111010011100011100", "01000010001100011010", "00110110100110011001", "01000010100101110111", "00111101111100110100", "10111001101100101001", "01000110111100010101", "01010010100100110111", "01010110011101011001", "11000010011100110111", "01011110000101000101", "00111110110110100111", "11100110000100010111", "11000110100100011000",
		 "01001101111100001001", "11100010000100011000", "10101110001011101010", "01001011001100100111", "11100110000011100110", "10110110011101101001", "01001010010110000111", "01001010000100111101", "11001001110100111010", "10111110010100100101", "01001001110100000111", "01111110110011110111", "11000110001100101000", "01011010000101010111", "01011111010100010110", "11000010000110001011", "01001010111011111001", "11000101110100001000", "10110110110011110111", "01010010110101010111", "01001010001100011010", "01000110011101011001", "00111010011100011001", "01001010000100111000", "11000011001100001001", "10101110001110000111", "00110010110100001001", "11000110000101110110", "10111001111100101101", "10110010000101001100", "01000110101100101000", "11000010010101110111", "11000010011100011001", "00111110001100010101", "01010110010100010111", "11001010001100101000", "11001110111100000111", "00111010111100000111", "01000110000100101000", "01001110110100011010", "01000110000100010110", "10111101110100100101", "01001101101110001000", "11001010001100110111", "11001110110011110110", "11010110110100001011", "10111110000011100110", "01010110000110010111", "11000110011011100111", "00111101110101111000",
		 "01010010011100111000", "11001110000100000101", "11000010011100001000", "01010110010011110101", "01000110101101011000", "11000011010100100111", "00111110011100111100", "10111010010100101111", "01000010011100001101", "01001010000100010111", "00101001101100101011", "11011111010100101100", "01001010000100010110", "01001011011100111001", "11001110100011101001", "01000101111100101000", "11001110101101011001", "01000110100100000111", "11000010101100010111", "01010010011101010111", "01001110011101011001", "01011010000110011101", "11001110000101010100", "00110010010100101011", "11000110101011101001", "10110110010100011100", "10111101111101001111", "00101001111100001001", "11001110000100001001", "11000010101101000111", "10111110001101001000", "00111001110011101000", "11011010101101111010", "10110110000100111000", "10111101111100101010", "11001110000100001001", "00101010010100000111", "10111010000100001100", "00111010110110101010", "01000110000100001000", "11000111001100100110", "10111110000011101010", "10111110011100000111", "11011010110100101010", "10111110000101111001", "11000110001100010110", "01001101101100100110", "11001001110100001000", "11001110000100010111", "01001010110011101001",
		 "11000010000101101000", "10111011010011111000", "01001010111100001000", "01001010011111000111", "00111110110101111001", "11000110010100001001", "01000010100100101011", "11000010001100001000", "00110010100110011000", "11010110000011111000", "11101110011100111000", "11000110110101111000", "00110110000100001111", "00111110011101101100", "10110110100100001110", "11010110000101001001", "01001101110110000111", "11001010011100100101", "11000110111110001000", "11011010101100111001", "00110111001100100111", "11011110001101101001", "00111011001100000111", "11000010010100110110", "11001011111100101000", "11000011110100011001", "11001110111101001010", "11001110011101011001", "11010110110101010101", "11001110100100100110", "11100110110100001001", "11000110010101011000", "01000010000100010111", "01000110001011111000", "10111110010100011011", "11001011000101011001", "01011010000100111001", "01000010001011100110", "11000011000100101101", "11000110100100000100", "11001110110100011000", "10110110000011111001", "01010010011100111000", "11100010000110001000", "11001110010100100111", "10111010011100100110", "11011010100100011001", "11100010101100101011", "11001110100100111000", "11000010010101100111",
		 "01011010011100101111", "11001110010100110111", "10111110011101110110", "00111010010100111011", "11001010011101011000", "10110001110100000111", "00111110111100101000", "11010111001100001000", "10111110101100101001", "11001011110100011100", "11001110011100001000", "01000110100101000111", "11011111000100010110", "11000011001011111000", "01000110111101111010", "11000010010101000100", "00111010001100100110", "00111110100100010111", "01000001111011111001", "10111001110100001010", "11000110001101010111", "00110110000110100111", "01001110011100110110", "01010010010101001000", "10111110000101111010", "01000110011110010011", "10111010110101011000", "10111010000100000101", "01010001110100110110", "01000110110100001000", "10101101101100001001", "10111010011100101010", "00110010101100111001", "11001010101101101000", "00111010100110000111", "11001110011100110111", "01000010001100010111", "01011111000100101001", "10111010110100110110", "10111110001011110110", "11010110101101000110", "00110010001100010111", "00110010000100001000", "01011010011110011000", "11000110110011100111", "11000110010101011000", "00111010111011000111", "10111010010100111010", "11000010001011110110", "00111101110100010101", 
		 "01001110010101111001", "01010110111100100111", "10110110001100101000", "01000001101011111000", "10111010110101011010", "10100110001100000110", "00111001111101110011", "10111110001101101010", "00110010010101000111", "11000101110100100110", "01000110000100101000", "11000010000011110110", "10111001110100111000", "00111110101100110111", "01000010001011110111", "01101110010110101100", "11100110101100110110", "00111110100100111001", "00111011111100011000", "01010001100011011000", "11100010011011001001", "10111110011110001001", "00111010010011100101", "00111001101100000101", "01000101110011000101", "11000001100100100110", "01000110000100110100", "00110001011100011000", "00111001100100010110", "10101101110011101011", "01001010000100010101", "00110001100010100100", "10111101100111010110", "11001001111011100111", "10111110000101110110", "11010010000100010111", "00110001110101000101", "10111001111101010111", "01000011001110100110", "00110001100100000101", "00110101111110000110", "00111011001100001001", "00110110101011000101", "11000110111101001011", "00111110010011110110", "01001010101100001000", "00101010000101100111", "01001001110011110111", "00110001110111101000", "11000101111011101001",
		 "01011010001100010111", "11000110000100001001", "00110110001011101000", "01001110101100100111", "01000010011101011011", "00111101110100010100", "00111010010101000101", "00111110001100001000", "11100010011011100111", "10111001111011101000", "11000001110100010111", "00111001110100010111", "01000001000101000110", "10101101110100101001", "01010010010111000111", "01101010000101011000", "00110001100100100111", "01001110010101000111", "01001101111111011010", "10110101111101001011", "01000110011100110111", "01000110010011111010", "10110101100101010110", "10110101111101001000", "01000001110100010111", "11010010011011001000", "01000011001011100111", "11000110011110011000", "11010010011101011001", "11010110000110001000", "11001110001101000111", "10110010101100001100", "10110101110110000101", "11000110010011100111", "01001110111101101000", "10111001100100001000", "00110010011101010111", "01001010010100000101", "11000010100101010111", "10111011010011111000", "00101001110100111000", "10111110001100101000", "10111101101011100110", "10111110101100110111", "01001110100011110111", "01010010111010100111", "11000010011100000110", "11010010001100100111", "01001001110101010110", "10111111000011010110",
		 "01000001110100000110", "00101110100101010110", "00110001110011001000", "01010110100110000110", "10110101110010101000", "01001010010100011000", "00111010001100011001", "00110110000101001000", "01000010000100010101", "00111010000011100110", "11000110100100010100", "00111110011101010101", "01000010111100000110", "11001111001100000111", "10110101110100101001", "00111001111011001001", "11001001111011010111", "10111010100110101000", "10111110000011101100", "00111001111100001000", "11011010000100100111", "00111010001011110101", "00111110100100001010", "10101110101100001000", "01001110110100110110", "11000110001100010111", "00111110001100101000", "00110010010100010111", "00111110010011010110", "00101101011011100110", "01100010000100011010", "01000110000011111010", "00110010001100010110", "00111001101101100111", "10110101110011111000", "10111010000011101001", "10110010110011101000", "00110001111100000110", "11001110011100011000", "01010010111011111010", "01000110000100100110", "11000110101011110101", "00110010000100101010", "01010110001011100111", "00111010001011101000", "01010110100101110110", "00111010001011010110", "10111101110101100101", "00111010110100010011", "11001010000011100101",
		 "01000101111101101001", "00111010000011000111", "10101001010100001000", "10110001111101000110", "11000010000011011010", "10111101100101000111", "01010010101101110111", "10110010010011000110", "00110110011011100101", "01000001110011001000", "01000001111110010110", "01000001110100010111", "00110101101100000100", "01101101111100001001", "00111101101011001010", "10110010000100011010", "10111010011100111010", "11000010000100101010", "01001010001100000111", "11000110101011111010", "01001010110100110101", "11000010010011111000", "01000001111011010111", "11000010011011010110", "01011011010100000111", "10110001111011100111", "10110101110101011001", "10110101111100011001", "00111010110010100111", "10111010100101010101", "01001110001100110101", "10111110000011111000", "11001110101100111001", "01000110001100000101", "01000010000110111001", "10111001111100010110", "00110110110100100101", "01011010000011110111", "00110010000011011010", "11000110111100110110", "00111001110100010111", "00111110010100000111", "11010010011100001000", "10110110101110000100", "01000010011100111010", "01000001110100100110", "00111010000010100111", "11000010000100001001", "01011001110100000101", "00111110010100000110",
		 "11010011000011110111", "01000001101101000111", "11000101110100011000", "01000001100011000111", "00101101110101011001", "11010010010101010110", "01000010110011110110", "01000101111101111011", "10101010110100001000", "11100010000101000111", "10110110000100110111", "00111110010100111001", "11010010011101110111", "10111110001011110101", "11000001111011101000", "01000110100011001010", "00111010000100000110", "01001010110011100110", "11010110011011110111", "11001110111011110110", "10111110111100110100", "01011110001100000110", "10110110011100010111", "11000101010100101000", "00101101111011011000", "10101110111011101000", "10110110000100001000", "11001101111100010110", "01101010011100000111", "01001010001100011000", "11000010100110001001", "10110001110100111010", "10110101100011011000", "10110010001110000111", "00110001110100011000", "00111110101100000101", "10111010110101001000", "10100110001100101001", "11000110001100011000", "01011010110011011101", "00110010101011101001", "11001110001011111000", "00101001111100100111", "00111110010101000110", "10110010100100001101", "01001110011011111000", "00101110010011100111", "10110101111100111010", "00110010011010110100", "10111010001011111000",
		 "11000101111100011000", "01011010011100100110", "01000010100111001001", "10101001100100001000", "11001010100111100111", "10111011001100111101", "01000011110101001011", "10111110001101001000", "00110101110011100101", "11000101010010100111", "01000001110011110101", "00110110001011111000", "10101110110011100111", "01010101110101011010", "11001010110101110111", "11001110001101011001", "10110110000111101001", "11000101110011010100", "10110110001100111010", "01011010000100011000", "10111010010100110111", "10101111010100010110", "01000010100011000110", "11000101100011010111", "00111110011100010111", "11000110000100101000", "10111110001011111001", "10111101101100100110", "01001001111100001010", "01000110011100011001", "00111010101100101001", "10111110001101010110", "11101010100100010110", "11000110110101001111", "10101110001011100111", "01000010001011111001", "01001101110100011000", "01000001111100100101", "01001110011100110111", "01010010010100010101", "10110110001100111010", "10101110001011100111", "11010110110100101000", "00111111011011010101", "00110001110011111010", "01001110001011110101", "10110011001101011000", "00111110000100001000", "00110010000101000110", "11010001110100001000",
		 "00111110011100000110", "00111010011101110100", "10111010000101011001", "00111101100100011101", "11010010011011110110", "00101001101011100110", "00111110100011100110", "01111010001100001001", "01100101101100001001", "11000101101011101010", "10111010111100001000", "10111010000010101001", "10110101101101111010", "01000001111100000111", "10111110110101000111", "01111110001011110110", "10110010100100010111", "00110010000011110101", "10110101101100001000", "00101001111011000111", "00111001101101111110", "00110001111100011000", "11010101110011010110", "01010011000100110110", "00111110100011110101", "01000110000100010110", "10110110111100010101", "01100010000110010111", "10110110010011101000", "01001010010011011000", "01011110010100000110", "00111010011100110110", "10110010000100110111", "00111001101100011001", "01000110001110010110", "11000101100111010101", "01010001110011000101", "01110001101101011001", "01000110011101010101", "10110101110100001001", "01010010101100100110", "00111010000100110101", "11000010010011101000", "11001001110100010111", "01000010000100010110", "11000001111011111001", "10101111010100011011", "11000101100100111000", "01000010110011101000", "00110110010100010111",
		 "01010110010100011000", "00100001111100100110", "10100001101011011000", "11000101110100101001", "10111110001011100111", "10101101100100011001", "11001110000100010101", "10111110001100111000", "11000011110100000110", "00101010000011100111", "10110110011100000111", "01000010010100000011", "10110010000011100110", "11010010111100001010", "01000101111011000111", "11000011110011100110", "00110110011011100110", "10110010100100010100", "11001110001011110100", "01000010000100000111", "00111110101011111010", "10101001110011110110", "01001101110100010111", "10101110000011110111", "11001101110011011000", "01001010110100000100", "00111110001100010101", "00110010100101000110", "00111010001011100100", "10100001111011101000", "01001001111101011001", "01001111000100100011", "01000011111100011000", "01000010111011110101", "11000110010100100111", "00011010010011000110", "00111101110101110100", "01011110110011100110", "10110010001100000011", "10111110001100010111", "00011001110101000110", "01000110011100010011", "00101101001011000110", "00101010010100001001", "11010010100011111001", "00011111011101000100", "11010001111100010110", "01010110000100010111", "00100111000011111000", "01001110011011111001",
		 "11000110000110010110", "00111010011011001000", "11001110001100110110", "10110110101100010111", "01000010111011100101", "11000010100011010110", "00110010000011010101", "00100010000011000111", "10110110010100110110", "11000010010011010110", "00110110001101010011", "00110010011101100111", "11001001010100110100", "11010001111011111000", "00111010000101110110", "01000010010100010110", "10111101010101001001", "10111110000101010100", "00110101100100001000", "10101101100100011001", "01000110100100010110", "00110001110011101010", "10111010011011000111", "10101001100100101010", "00100001111100110110", "11001110101011010110", "00111110000011110110", "11001110000100011000", "00111010011100100100", "00111001111011110111", "10100101111100010110", "10111110001100111011", "10110001110101010101", "01010110001101111000", "10110010110100000011", "00101010010011100100", "10110010000100000101", "10110110010011100110", "01010110011100010100", "10101001111011001000", "10101110001100110100", "00100101111011100111", "10110101111011110110", "01000110010100000111", "11100101111101110111", "01001110001100010111", "10100010000100011010", "00110010000011000101", "11001110001100100111", "11001110000100010011",
		 "10111110011100000111", "01001101111100110110", "00110010011100000110", "10110010011100100110", "10111101111100001000", "01000101111011010110", "10110010000101110111", "10111110110101010101", "11000110111100110011", "10111010000011010100", "00110010011100100010", "11000110100100100111", "01001010001101001000", "10110110111100011110", "11010001110011101100", "00111010011100010101", "10111110001100001011", "00111101111011101001", "10100110001011011000", "10101001010100000111", "10110101101011010101", "01000010001100000110", "00101010000100000111", "11010010101011010111", "01000110100011110011", "01001010100100010111", "00101001101100101000", "11000101101100000101", "10111110000110010101", "10110101000111101001", "11001010001100110101", "01001001110011111010", "11000110100100111000", "10111010000100010101", "00111110011011000101", "10101010011101100110", "10111101110010101001", "00101010001100010111", "01000010001101010111", "00110110010100110101", "01001010010101000101", "10110001100101001000", "00110110101101000100", "00110001110101010111", "00110010011100010111", "10100110010100110111", "11010110001011100110", "11001010001011100011", "11001110110011110101", "00111001110100110110",
		 "01000011000101011000", "10011101100100101001", "10110110010011110110", "00100011001011000100", "01001110010011111000", "00111010001100000101", "01010010010100010111", "10111010010011111000", "01000110011100100111", "00101110101101000100", "01000001111011100100", "01001110000111000101", "00101110011100110101", "11100101110100101000", "00110010011011110110", "01001001111101001000", "10111110011110001000", "00101010111011011001", "00100111011110100111", "00110110100100100101", "00111011100011100110", "11000001111100101000", "00111010001101110110", "11001110011011100111", "10110101111100010110", "00101110011011100111", "10111010000011001000", "01000110010011110110", "00101101110011000110", "10110010000011010100", "10110110101100010110", "10111110000011101001", "10100110000100010110", "01010010011101110100", "10110010000011100011", "00111001111011010111", "10111001110101010111", "10111010010100010110", "10111101100101000110", "00111110011100101010", "00110110100011010100", "01000110100100000111", "10100101110011110110", "11000101111100100111", "01001010001100000101", "00110001111011110011", "10110110010010100110", "10110101111100101001", "10110101010011101001", "01011110101010100111",
		 "11010010101011111000", "01011010010011000101", "00101001111011000111", "01001101110100100101", "10111010010100110110", "10111001101101010110", "11000001110011100101", "00101110011100011000", "10110011011011100111", "10101101110100101111", "00111111000011001000", "10110110011011000101", "00111110010100010111", "11000110101100011000", "00110010000100101001", "11001110010011110101", "00101010111100011011", "00101010011101110111", "11010010001100001000", "10110010110100110111", "11001110010101000110", "11001001111100010101", "11000110101011110100", "00100001011100100111", "00111110011100101001", "10100110101101100111", "00101110100100101100", "00111001010100111000", "10101110000101010101", "11010010111100000111", "00110010001011101010", "11011010000101011000", "10110110000101111000", "10110001110101101001", "01000010011101010101", "10111001111100000110", "00100010100101011010", "10110001101101001000", "10101101111011010110", "11011010010100010110", "00111011001101011001", "00111001111100000110", "00101001111100100100", "11000001111100001001", "01001001111101111011", "11001010000011111001", "00111010111100100100", "01001010010011111011", "11001101111101000101", "00101010001101011001",
		 "00111110010111001010", "00101010000100011001", "11010010001011111001", "01000110011011011110", "10110001010011110111", "00101001110101100101", "11100101100011111000", "11001010000101011101", "00011101111011110101", "11010001110010000110", "00110001110110001011", "11010010001011100111", "10110010000101011010", "01000110101110101010", "10110110000011110110", "10101110101100111100", "10111001111100000100", "10111101101101001000", "11001110000100010110", "10111010000011000110", "00110110011100111000", "01001010001011110110", "01010010000011100101", "10110101100011100110", "10111110100110110110", "00111110000100011001", "10111110000100101000", "10100110101101100110", "11001010011110010011", "11000110011100000011", "11011010001011100110", "10110110000100001000", "11000010010100010101", "11010010001100101101", "11001010000011111001", "01111010100111110110", "00111011000100010110", "00111001100100100101", "10110110011011110110", "10101001110101000101", "01111010010101001010", "00100111011011111000", "10111101111100010110", "00101001111100000101", "10101010001100110100", "00110010001101000100", "11010101101011101001", "00111110010011100101", "01011110000100011001", "00100010011110000011",
		 "01001111001110010101", "11000110101100110101", "01001110011101100101", "10110101100100000100", "00111110010100110101", "10110010111011000101", "00111101010100000101", "10110110110100011000", "10111001111100000110", "10101010000101101001", "10100011000011001001", "10111001110101011001", "00110110001011010111", "10100010101110011101", "11000101111100110110", "00111110101011110100", "01001010000011101000", "10110001110011110101", "10110101111100000110", "00100101110011001000", "11010010000011100110", "01000111001100000110", "00101010000011100101", "00100001101011100111"); 
		weight_ROM(9) <= (
		 "10110101100100011010", "01000110001101001001", "00110001011100011001", "01000110001100000111", "01010101111101011010", "10101101101101001010", "10111110000011100110", "00100010001100000111", "01000010110011101000", "10110010000100010111", "10111010001100101010", "11001110000100000101", "10110010010101010101", "10111101111100111000", "00111010010100111001", "11000010000100100111", "10110110010100010101", "00111010000100010110", "11000110001100010111", "01010110010011110101", "11000110001011110101", "00100101101100000110", "01111110001101001001", "00101110111100100111", "11100010010011010011", "00110010011100001000", "11001010100100110101", "11010110010100001100", "00111010000100010101", "10111010010011101000", "11000010100100001001", "11010110000011010101", "01000010001100100111", "10111110000100110101", "01011010000110011010", "10101111000011101000", "10101101000111000101", "11001010001011111010", "00111110001100000100", "01000110111101011001", "10101110010100001000", "10111110001100010110", "00100001111011001000", "00101110010100010110", "01010110011101010111", "10100101110011100101", "01001110001011100111", "11010010011101011010", "00100110100011111010", "01000110001011101000",
		 "11001010010100010111", "10111110001101001001", "11001001111101011010", "10110111001101100101", "01000110000100110111", "01000111001011110110", "00111111010011000110", "10111111010100010100", "11001001110100110110", "10111001110011001000", "10110010001110010110", "01001011001011111001", "11001110001101110101", "00110001110011101011", "11001011000100111000", "01100001111101010110", "11010001000011101000", "10100011001100110100", "00110101111100001000", "10110010010110111000", "00111010000100101000", "00101010110011100101", "01000010100101000111", "10101101111101101101", "01000110000111110100", "00110010010101000110", "10111110011011110110", "11010110010011101011", "10110110000100100101", "11001110000101010111", "10101110010100111000", "11001010100100001001", "10101010111011101001", "00111011010110101000", "10111010101100010101", "00111110111011100111", "00110111000011100110", "10111001110100101010", "10111110000110100100", "01001001100011110111", "00110001111101011010", "00111011010100010110", "01000111101011011000", "11001110001100010110", "01001110010100000101", "10101010000011010111", "10110010011100011010", "11001010001010100111", "00111010011100011001", "11000110000100110111",
		 "00101110001100100011", "01000001110101000111", "11001010000100111010", "10101010001101010111", "10111101111100001001", "11001010011100110111", "01010010100100010110", "00110110000011011001", "11010010001100010100", "01000110010011100101", "01001001111100100011", "01001010011100101001", "11100010001011101010", "10110110100100101010", "11101001110100101010", "01000101111100000111", "11010110111100101001", "10110110110101101000", "10100010000011011000", "11001010001100001010", "10111110000011100111", "00111010001011010111", "10110101110100011000", "10111110000100101001", "01001110000100010100", "01000010001101000111", "10111010001101001011", "10111101111100010101", "00100001110100100101", "10101101100100011001", "10111101110101000110", "00111010000011110111", "01000101111101111000", "10110001110100010101", "10101110001011110011", "00111010001101000111", "10100001110100011010", "00110010010100100111", "00101001101011100111", "11010010000111100101", "01001010000100000110", "01000001010100000100", "10111011001100000111", "01001010101101000101", "11010010111011110110", "00111110010100110101", "10110110000011111100", "11011010100100110110", "11000110001011110100", "00111010111011100111",
		 "11000110011100110110", "00110001111101100111", "00101110000100101001", "00110110000101000110", "01000110010011100101", "10111110001011010100", "01000010000100011000", "00100110010100100111", "01001101101100010111", "11001010010100000100", "01000110001110010101", "01000010010101010111", "01011001100011010100", "11011110010100101000", "01000010111100010111", "10101010011100011001", "01010110100011111000", "10111101010011010110", "01000010000100100100", "00111010100101000101", "11010011000101101000", "10111110001100011001", "01000010010111110101", "11010001110100000111", "11011010001011101101", "10111010011101111010", "10110110000011011001", "10110010001101110100", "01000010000100000101", "00101001111011000111", "10101010000100010110", "01010011001011110111", "10011110011100101000", "00111110011101010110", "01011010100100010111", "11001010011100010110", "11000001101100101000", "00110110010011010111", "00110001111100100110", "01000010010011110110", "11000110000011000101", "01000010001101000011", "01010101110101111010", "11010110100100111100", "01001010000011011010", "01000110011100010100", "10101110100010110110", "10110010011100111010", "11000110010100000101", "11001010001100110101",
		 "00111001111011100101", "11010010100100000111", "10111110000100101001", "01001110010011110111", "11000010011100001001", "00111010011100100110", "11010010000101101000", "00111010011100001000", "10111001111100011100", "10111010000110001001", "00100001010101101100", "10101110010100010110", "11001010011100010110", "01000110011011111000", "10111010000100101001", "01000001100011110111", "10101110010101001010", "00110001110011001100", "11001010001011100101", "00111110100011101001", "01111101110100010111", "10111001111011100111", "11000010001101010010", "00110110111011101100", "10110010011100110101", "10011010000100110101", "10101101101100001001", "00100010001101001001", "11000101110011100110", "11010010010100110111", "01000110011011000110", "01010010000101011011", "10110110010101011101", "10111110100100101001", "10111101110011110111", "00111010011100100110", "00101010000011111001", "10101010101100111001", "11000010001011010111", "00110010001101010110", "00101010111100000111", "01001011000100110110", "00100001001100100100", "01001001110100111000", "01010110000011111001", "11000010010101001000", "00111110000100100110", "10101101111100001011", "11010011011011100101", "01010010000100011000",
		 "10111010100100011001", "11000010101100011001", "10111010010100001000", "01101101110011100110", "10110110001101011000", "00111001101100001000", "01100110100100011001", "11001010001100111001", "00100101111100010101", "01001101010100011000", "11010010011100001011", "01001010010100110101", "01000010110011001100", "11000110011011100111", "10111101010100110100", "00111010010101001010", "00110110011100010100", "11100101110011110011", "10111010010100011000", "11000110100011100111", "00110110000100100110", "10111110011100110101", "11001101111100100111", "10111101100011010111", "00110110100100010100", "10100110000101011010", "00111001111100111011", "00111011010100000111", "11010010001100010101", "10110110000100100011", "01000011000111100101", "10110101111101001011", "01000110101100010101", "11001010011100111001", "10110110010100011010", "11001010001101010111", "11010010000100110111", "00110110010100001000", "01000010000100010101", "10011010011101111000", "01010111101100001011", "10110010000100101000", "11000010001100100101", "00111110100100100110", "00100010000011000110", "10101110010100100110", "01010110001011101010", "11000010001100111010", "11001010101100000111", "10111110100100111000",
		 "01000010011011100111", "01001110001100110101", "00111010111100100110", "01010101101101110111", "00110010101110001000", "00110110100100010110", "11000010111010100110", "00110010100101001001", "11001111000100000101", "10111101010100111000", "10100001110100011010", "10111101110011100111", "00110110001100001001", "10110001101100000111", "11101101110110011001", "00111010001011000100", "01100011011100100101", "00111010100011000101", "10101001101011101000", "10101001101100011000", "00111110000100001000", "00101110011100100111", "01001011000100010110", "01011001110100000100", "01000110010100100111", "11000110110100010011", "00111110011100110111", "01100010000011110101", "00101001100110010101", "01100010000100100101", "10110011000101001001", "10110010111100001010", "00101110110100101001", "01010110001100001000", "11000010000101010111", "01000111000101110110", "10110001110110000111", "11010010001101001111", "11010110101100010110", "00110001111011010110", "10110010001100101001", "00111110100100110111", "00110110110100001001", "11001110001011101001", "11011010000011110110", "10110010010101111101", "00100010001100100110", "10110110000100101000", "00101010001100110101", "00111101110100010101",
		 "01110110011100001000", "00101101011011001001", "00101001010011100111", "01001011011011110111", "10110001110011101000", "10110101101110001001", "01011001111101110100", "00101110010100100111", "01000110000100110111", "00100110000101001001", "10101001110100001000", "00110010001100110100", "00110001111011000111", "01001010001101100111", "11000010101101010110", "11001010100011110110", "00110001111011101000", "01000101111101000110", "01001001110100010101", "01001011010010110110", "10111101111100111001", "00110101101100011000", "01010010010100010111", "10110010001100011010", "01000101111100110101", "11001010011100110110", "11001010001100011000", "01011101110100110110", "10111010011100010101", "10101101101101111000", "11001010001100100111", "11011110001010100101", "11000001110101111001", "00110001110100111000", "01010110001101101000", "00100010101010100110", "11000001011100010110", "01010001110100000101", "11000110011101000100", "11001110110100110110", "10101010001100001001", "11001010111101000111", "00100001101100100111", "10101101110100110110", "01001110001100110111", "00101010100101010110", "01000001111100000100", "00111110001101110111", "00110011001100100111", "10101101101100001011",
		 "01001110010100111000", "10110010001110001001", "00111001010100010101", "11011110010100000110", "00110110011101110011", "00111010100100011000", "00100001110011100110", "10101010110100000111", "10111001110100100111", "10111110011101101011", "10101010100011100100", "01111111000100001000", "00110010001011100100", "01000001110100001001", "01001110011100100101", "00110011101101010101", "00110010001100101010", "01010110011100110101", "00101101100100011000", "00110010001011010110", "11001010000100110100", "00101010000100100100", "10111101110100001010", "00110101111100001000", "01001010010011100101", "01011001110100010110", "00110011000100111001", "11001111100100110110", "01001001110100111010", "00111011011100011000", "10101101101100101000", "10111101111101010111", "01010110111011100110", "11001110000100110110", "00111110000110000101", "00111110001010110111", "01000110010101010110", "00111110011100010111", "00111011000110010101", "00111001110011011000", "10100001100100101000", "10110001111101100110", "01100010101100010111", "01001110000100110101", "11010010000100110101", "01001001101011011001", "00110001110100101000", "11000011000100100100", "01011010010011111000", "10111001110100100111",
		 "00111110011100100100", "00111001111101110101", "00101001111101000110", "11000001111011110100", "10101110110010101011", "00111010000100100110", "00101010100101000110", "00101110000100000100", "01001010010011010100", "00111101110011100100", "11010001111011100111", "01000010001011110110", "11000010011011110110", "11000010001101101001", "11000101111100001001", "01010010011100010110", "11011110111010100100", "10110010111101001010", "10100011010100011000", "00110101110011001000", "00110001111011101001", "01001110011100110101", "00101010100100100101", "00111111010011101001", "00101010000011110101", "11010110000011000100", "10110101000101000111", "11010110011011110100", "10110110000011110101", "10110101100101011010", "10111110011100001100", "01000001100100110110", "01001010000101010111", "10100110000100000111", "00101101001011010101", "00110101100011110110", "10111001111110011000", "01001010001101110100", "00101010001100000101", "01000010000100100101", "01000001010011110011", "00110001000100101001", "11010110000011100101", "10111101011011101000", "01000110111100110111", "00100010011101101000", "00110110000100000010", "11001001111011010111", "11000010010100010011", "10110101110110110111",
		 "00111110001110010111", "00111001101100100101", "10111011010100001011", "00111111010011010111", "00111001100100101010", "10111101110011110101", "01001010000011110110", "00110001111011100111", "11010010101011100110", "01001011000101000100", "01010110010011110101", "01000110111101010100", "11001010001010100100", "11011010001100011001", "11000110000100010011", "10110010100100000111", "10111010000110100101", "10011101100100011001", "10101010010011110101", "00111101100110100110", "01010010011100010101", "11000001110101001001", "01001111010100111001", "10111010010100111001", "10101110011100010111", "00110110001011101001", "00101101100010101011", "10101110000101010110", "01001010001011000111", "01001001111010110110", "01000010100100100110", "11000101110011100111", "10011110000100001000", "10111010001011000110", "11000010000011001000", "11011010111100111010", "01010010010100101010", "10111110010100111000", "01001010110100100110", "01000010001011110101", "01011110010011000100", "01011111100100100101", "11000110001011110111", "11001010001100010100", "01011110111010100101", "00100101111011000100", "10100110010010100100", "01000110001101001001", "10101101100100001000", "00111110001100110101",
		 "11000010000100110111", "11001110010100100100", "10101001110100111001", "01001101111011010100", "11011110111100110111", "00111001111100000100", "00111011100011100111", "01001110101100111001", "00101110111010100110", "11000010101100001001", "10110001100100011001", "11000110011100010100", "10111101110100110101", "01001010011101011001", "11000010010110010110", "01010110100010100101", "00100010001100100111", "00111010001100000101", "00111010111100010110", "01010110111101111001", "00111010001110011000", "11000010000100100111", "00111010000100010110", "00110101111011100111", "10110001111100010100", "10101010001101010110", "10011101100011101011", "00101001101011110111", "11001110101100100110", "01010110001100110111", "10111001111100100101", "11010110001100011001", "10101010001100011000", "01010010110100101101", "00101110010011010101", "10110110101011010101", "00110001110100100111", "10101110100100111010", "00101001110010100101", "00110010000011000110", "10110001111011100100", "01000010010100110111", "11000000110101100110", "10110010110101000110", "11010101111100111000", "11011110100011111000", "00110101101011100101", "10101010011100001000", "10111110111100000100", "11010010100100001000",
		 "01001010000100011000", "01000101100100011000", "11000010001100011001", "00110110010100010101", "10111101100100010111", "10101110111101010111", "01010010011110110111", "11101110110100001011", "00100001011011100011", "00101010011101011001", "11000001110101111000", "00101011011011110111", "10110010100011111001", "01000110010100010111", "00110101110011111100", "10110110110100111000", "00110011000100100110", "00101110111100110101", "11000010111011011010", "10110010001101011000", "00111010000100100100", "11000001110100010011", "00101110000110000111", "00111101100011010011", "10110010000110110011", "10101001111011111010", "11001110100100101000", "10110101011011110101", "01001011011100010101", "10110010110100001000", "01000101111100100110", "10111101111011100111", "11000101111100100111", "10111011000100110111", "11000110100011000100", "01000101111100010111", "01100101110100010111", "00111010000100000110", "10111011001100010111", "10101010011100100100", "01001010111100001010", "10100110011100101010", "10110001101100000110", "01000010001100000111", "00101110000100000101", "00100101111100000100", "00110110001100111001", "10101001111100100101", "10111010001101010110", "11000001110011110110",
		 "01000110000100110101", "00111110001100010100", "10101010001101100110", "10110101011100100110", "01001110000011110010", "10011010001101110111", "00111001110010100100", "10111110000101011001", "10110101111011001001", "10101101101100011000", "00101111101011100110", "11000110001011001000", "10111010010100011000", "01000001110111000110", "10111110001100100111", "10110110011011100110", "00110001110011100100", "10110110100010100111", "00110101100101000111", "00111010001100000111", "11010111001100111000", "10110010011011111010", "00111001110011010100", "11000001100101100110", "01001010011100100101", "01110001110101010011", "11010010000100110111", "10111001111100010110", "11001101100011010100", "00101010000100010100", "10111001111011100111", "10111101110011111100", "00110010011100100100", "01000110011100000111", "01001010001101001010", "01001001110101010101", "10111110000110110110", "11000110000101011010", "01000010001100110101", "00110001111100000101", "00110101111011110011", "11010111000101110111", "10110001110011001000", "01001010011100111000", "01001110000011000100", "10100110000011001001", "00101110000101010111", "01100010100101000101", "00111010011101010011", "11000010010101010101", 
		 "11011110011100111001", "10111110000100101000", "10101001111011011000", "01100110010100100101", "11001110000101011001", "10101101101100001010", "00111110000011100101", "10111111001100101001", "11010110100100001001", "01001001111100100111", "10101101111100101001", "00111010011011100110", "00110010001100100101", "11001010111101001000", "00111110111100000111", "00111110000011110110", "01000010111101111010", "01000010010101011000", "01000110010100010100", "01000010100111110101", "01001010001100010111", "10100111011100011110", "11010011100011111000", "01000110000101000111", "00111101010100010110", "00110101111011111000", "11001110110100010101", "11000110000101111000", "11000001110100000110", "10101110000100011001", "01000001111100011000", "10111010000011010101", "01001110001100100110", "00111010011101011000", "00111110000101001101", "00100110010011110110", "00110101010100110111", "01001010000100000111", "10101001100100100011", "01010110111100010110", "00110110110110000111", "11000101111101000111", "00111101101100001000", "00111010101100000110", "01010110011100111000", "00110010000100110110", "01011110100100010101", "01001101110100010111", "00110011000011110111", "10110010000100011110",
		 "01001010001110010111", "11000110100100011000", "01000001100100100110", "11000010010110010101", "01000110001100100101", "01000010011100000111", "00110110011100110101", "00110011111100000101", "11000010011100010110", "10101001110100100111", "01000111001100110101", "00110010011100000111", "01010001010101010111", "01001001110011101000", "11001110100101010101", "11010110001100110110", "00101101010100001010", "11000010101101010100", "00100101110100001000", "10101101111011010111", "01000111101100010110", "00111010001101010110", "11000010101110110111", "10101001110011111001", "00110010001100110111", "01001111000101001000", "01000110000011100110", "11010010101011101001", "11110001110100110111", "00110010001011111001", "10110001111101001100", "10111011000101111000", "10101010100101100110", "00111010010100110111", "00101011011100000100", "00110010111011100110", "11000011000011100100", "11000010100100100110", "00111010010100110100", "00100110010010111000", "10011010110111011100", "10100110011101000101", "10111101111101110110", "00111010110100100110", "11001010011100011000", "01011010001011000101", "10111011110100010111", "11001010010011000011", "11011110001100011101", "00111110010100110100",
		 "00110110001011011001", "11000110000101100100", "11000101111101000111", "10101010001100110110", "00111010101100101001", "11000110110100001010", "01100101110100000101", "10110010001100110101", "01001001110101011000", "10110010001100110101", "01000001111100000110", "01001010000100100101", "01100001110101010101", "00110001111100000111", "11000110010100111000", "01000010011100000101", "01000010110100010111", "11001010010100101000", "00111010000011011110", "10111101110100101001", "11000110011011100111", "11000110001100000110", "00110111001100100110", "10111110001101101001", "10110010110101011001", "01000110011011110111", "00101111000110011000", "00111001001100100100", "10111111001011100110", "11000101101100001000", "11001101110100010110", "11000001110100101001", "01000110100100001010", "10111010000100010110", "00111001011101100101", "01000110111110101001", "10110110010011101001", "00111011101100110111", "11001001101110000110", "11001110101011110100", "11001010001100100011", "01010001101100110111", "00101110010011100101", "01000001110100000111", "11010110101101000101", "10111110000110001000", "00111001110100010110", "10110010001101010110", "00110010101100010101", "00110010010100100110",
		 "10111110011100110110", "10110110000101000101", "10110110010101001001", "11000110011011010111", "00111110100100000110", "00110001111100000110", "01001111001101110110", "00101010100011111110", "01000010001110011000", "00110010010101000100", "01000101011100000111", "00111010101100000100", "01010001101011110101", "11001101110101001000", "00111010001100110100", "10110010100101001000", "01010010000011100111", "00110001001100000111", "00101011001011100110", "10110010110011100100", "11010010001100010110", "10101110000100011110", "00111001110100010101", "01001101111100101011", "10111110100111010111", "00101010010101101001", "10110110001011101001", "10111110100011000101", "01010110000011010110", "10110001010011011000", "11001110011101010111", "11100110000011110111", "00101001101100000111", "00111001110011110110", "00110110100011100110", "10111010000101100101", "01010001111100110110", "11000010000100010100", "10110101100101001010", "11001101111011110100", "00101010100010110110", "00111010000100010011", "11001101101011111000", "11001010010011100100", "01001010100100000110", "10101010101101100110", "00101110010011010101", "10111110011100010111", "10111010101100110101", "11010101111100100100",
		 "01011010001100100111", "11001011000011100011", "10111010101100011000", "11011101111100000111", "10110110100100110110", "10110010000011111000", "11000010000011101000", "00100110100101111000", "10011010100110000111", "10111010101111001001", "00101001111101001001", "00101010001100000110", "10111010001011010110", "11011011111100011000", "10110110011100100111", "00110010001101100111", "10100010000100010111", "01010110100100110100", "01010110000110011000", "01001110100110001011", "00110010011110101010", "11010010001100111010", "01000110011100110100", "00100110001100100111", "11001001111011010101", "10011010101011100110", "00100101111110011011", "11010101101101000111", "11000110000110010111", "11010110001100110110", "11001010000100000111", "00111010000100101000", "10110110001101001101", "10110010001100001000", "11000101110011000110", "01011110011100010101", "00101110011011100111", "01010001110101000111", "11001110000100100111", "11100111101100010110", "00101011001011000011", "01001010010100001100", "00101001011011100101", "01100001110100001000", "01000110011100001001", "01000111000100110111", "10110101100100011011", "00101001110100000111", "00101010101100001000", "00011010000101011011",
		 "11001111000011101011", "10101001101100111001", "01001110101011111110", "00110110001100101101", "00110101110011001011", "10110110111100110110", "01000010000100101101", "10111010001100111011", "00101101101100101011", "01000101110011000110", "00111110011100001000", "10101001110100010111", "00101110010100001000", "01000010101101100110", "10101101110110010101", "10111010100101011000", "10111110010110010110", "00110011000100100101", "01001010101100000110", "10110010010100010100", "01110011110011110110", "11011001111011100101", "11000110010101000100", "01000101101100100110", "01001110000101110100", "10111110011101101010", "11000010010101011001", "10101110000100110110", "00111110100100110110", "00110010010100100101", "11000110010100111000", "10110001111100010101", "11000010011011110101", "10111010101110001011", "10101110010011100111", "00110010011100000111", "01000110011100110110", "10101010011101000111", "10110110110100000110", "01000001111100100101", "10111110100100111001", "10101001111101011010", "01011010000100001001", "00101001101101010111", "10110110000100010101", "10100110010101100011", "00111101111011111001", "00100110101100100110", "01101110001100111000", "01000110011100100101",
		 "11001010010011110101", "00111111001100100110", "00111110001011010111", "00100001101100100100", "10111010111101010110", "10111010001100000111", "01001001111011100101", "11001010000100001000", "00110010001100000111", "10110101010011110111", "10100111000110000110", "10110110110101011000", "00110010001100000111", "10100010111101011001", "00111010010100011000", "10110110011100010101", "01001110010011110110", "10111010000011100111", "00100110010101101000", "00101001110100111010", "11101110010100000111", "00110110001011000110", "00100010100010100100", "01000110000100001010"); 
		weight_ROM(10) <= (
		 "11001110000101101000", "01000110100101001001", "10111101111100100111", "01000010001100010111", "11010010001110011001", "10101110000100101000", "00111010110011110101", "01011010111100101000", "00110010011101001010", "11000101011100100111", "00110001110100000111", "01010110011011100111", "11000010010101101111", "01001110011100001000", "00111010001100110111", "01000110001100101010", "11001110101011110110", "11001010100100101000", "00110110110100010111", "01010010000011010101", "11001001111011111001", "11010101110101011000", "01001010100011100111", "00110001101100010111", "11011110000011000110", "10111111100100000111", "10111110101101110100", "00111001101011110111", "00110010001101011000", "10111110110110101100", "01000110000100110101", "00110010010011100111", "10111101110101011000", "01010010001100010111", "11001110001110110110", "10111110001100111010", "11010001101110100110", "01001110101100111000", "00111010001100100101", "00111010010011100100", "00100101111101001001", "00110011000100001001", "00111101101100000110", "10111010010100001010", "01110111001100010101", "00111010001100001000", "00110001111100001000", "00111010000011111001", "00101010010100111011", "11000110111011111001",
		 "11010110000100011010", "10111101101101011001", "00111101100101101001", "11001110101011100110", "01001001100100001000", "01000011000011110101", "00110011000011101000", "01000001111110100110", "01001010001100011000", "01000001111011101000", "10111010010100111000", "01001010100111011100", "01001001100011100111", "10101010011100111001", "11000010000011110111", "11000110010111111010", "00101001111100000110", "11001110010100001111", "00110110000101001000", "11011010101100111100", "01001110101100110111", "01000010000100000110", "11000111000110010110", "10110101110101001001", "00111001110100001000", "01001010011011100111", "11000010001011111000", "01010010010101010111", "11100110010101011000", "11011110111100111001", "01000010111100100110", "01011010001011111110", "10110101101011100111", "11000011110011000110", "01000010001100010111", "01000010000011001000", "01000110001101011001", "11001110000011000110", "11000010101100010101", "11000010111100101000", "00110001110100001001", "01010110110100000110", "10110101101011100101", "11000111101100110111", "01010010000100010111", "01000001100011000111", "01111110100100011001", "00111110100100001000", "01000011010100010110", "11001111000100010110",
		 "01000010010100000100", "00110110000100010101", "00110001100011001000", "00111110001101000110", "10101101100010111000", "11000010100110011000", "11011001101100110111", "00110110010101010111", "00111010101100110110", "00110010000011100111", "11101010010100110110", "11000010000100110111", "01001110100101011100", "10111110101011000111", "10110101111100011000", "01000010011011110110", "01100010001011000111", "10110010000011001011", "11000110000011000110", "01000001101100001000", "01100110000100001010", "01000010001100110111", "01001010001100001010", "10101010011100001000", "01001110010011010110", "01010110101100011000", "00101110011110000111", "00110010000101011001", "01000010110011110110", "00110101011011000110", "01000110110100111000", "11100110010011111010", "00110010001101110111", "00110011011100111001", "10110101110011101001", "10111010100100000111", "10101110010100100111", "00110010001100100111", "11000010011011101000", "00111010001101100111", "01000101101101000111", "01001101111100110101", "00110001110100001001", "00111010101011000111", "01000010011100001001", "11010001111011110111", "00111010101010110111", "01011101111100000101", "11001001110011010100", "11001010000011000110",
		 "01011010101011111010", "00111101110100000111", "10101001110011101000", "10101010011101011010", "01000010000100001001", "11000110000100101000", "11000010101100010111", "10111110000011100111", "00111110001100111011", "11000001110011110110", "01010010011100000111", "00111010000100001010", "01000101011011100111", "10111010001011110111", "00111110101011110111", "10101110010100011001", "10110101110101001011", "11001110011100001001", "01000110101011001000", "11001010001110011001", "01100010100100010101", "10110101111110010111", "01000010001011110110", "11001110001011101011", "01000010000100110111", "01000001101100000110", "01010111011100011000", "11000110001100010111", "00110010000011000110", "10101110110101111000", "01010010100011111000", "11001110010011111011", "11101010010100111010", "11100101101100010110", "00111010100100001001", "11000001111101011000", "11001001110101011010", "11000010100011011001", "00110010001100100111", "01101111000110010110", "00111110110011110111", "00110110101110011001", "11000010001100101001", "10101010001011100111", "11000110011100111001", "00110010010100001000", "00111010010011011000", "11000010001100000111", "01000001111011100100", "01000010001100100111",
		 "10111101100100010111", "00111010010100001000", "10111101110100001011", "01001010000011101011", "00110110001011111000", "11000010010011110110", "01000110010110111000", "00111010101101001000", "10101101111100001010", "01100110010100000111", "11000101110111001110", "01000101111011101010", "10110101110101110101", "11000110011011111000", "10111010001101101000", "11000101110011110111", "01010010001101001010", "00110010010011100111", "01000010111011101000", "11000010001100010111", "01001010000100010110", "01011110011011010111", "11010010001100010101", "00110101110100111010", "00101111011010100101", "10100110001011101000", "10110101110011101000", "10111101101101110110", "11010010000101100101", "01001110101100110110", "10111010101011101010", "10110010101100101100", "10110101110011101001", "11000001110110011101", "00111001100100000110", "00110110011100000110", "10110001111100100111", "10101101111100111011", "10111110010100011001", "00111110000100010111", "00111110111100100110", "01001010110100010111", "00101001011011100110", "00111010001011000111", "11000010100100101010", "11001101110110011000", "00101110000011100111", "10111110001101000111", "00110010001011010101", "10101010011011010110",
		 "11001011000100011011", "00110001101100101000", "11001110101100101010", "10101001101110000111", "10111001110100100111", "10110010100011101000", "00111010010110111000", "10110010110100101000", "00110110000100000111", "01000101110011000111", "00111010000011110111", "01000010011100011000", "10111010000011101000", "01010010000011111000", "11011110001110111000", "11000101111101011001", "10111010001110011000", "11000110100011110110", "10110101111100110110", "01001010100011111000", "11000110000110000111", "10110111011101010110", "11011110000100011000", "11000010110011101000", "01011110001011101011", "11000110010100001000", "11000010101100101101", "11000101101011100111", "01000010100100111001", "11011110011011100111", "00111010001101101000", "11000110011110110110", "01000010000101011000", "11000010000100011000", "10110001100101000111", "00111010001011110110", "01001110011101111010", "01101010000011100111", "11000111011100010110", "00111110010100110110", "10111110001011110111", "10101110001101011001", "11001010101100011011", "00110001111011010111", "00110010000011100111", "11100110001100010101", "10101101111100011001", "01001010000011000101", "01001010000100101000", "01000010001100100111",
		 "11001010011101000110", "01000010001100010110", "01000010100100100111", "01000110000010100111", "01001001111100110111", "00110010001101100110", "01000101100100100110", "10111110011100011000", "10111101100011000111", "10111101111010101000", "10110110000011111001", "10101010001011100111", "10111011110011110111", "01000001111100000110", "10111010011101001000", "01110110101011010101", "11000010110011111000", "00111010000100010111", "00110010011100100111", "00101001101011100101", "00111001101100000110", "00110010001100110111", "11001101110011110110", "01000010011100010110", "10111110000101110110", "00110110010011000111", "10111110000110110110", "11001010000100110111", "11001101100011100111", "01000010000100010111", "11000010010011100111", "00110111011011111000", "10110111010100110111", "00111011101100010111", "01000110010011110110", "01010101110100110111", "10111001110011000101", "01000010011100011000", "01000110011101100111", "10110110011100111010", "01010010001101001000", "00111101110100010110", "11001001010011100110", "01000001111101010110", "01000011110011110110", "01001001101100001100", "10110010001011101001", "10111110010101111000", "11010110001100100101", "00111101110100010101", 
		 "11000101111110001101", "11000010000100001010", "01011110101100001111", "01010011110100101010", "11010110101110010111", "01001001111100101000", "01011110100110110110", "11000010010011101100", "00110010010100111010", "00110110000100111001", "01001101111101101010", "11001110101101000110", "01001010001101010110", "11000010100100001000", "11001010001100010111", "11101010001100111000", "01011110101100101000", "11001110100100101001", "01011111000100010101", "00111010100110100111", "11001110011100001000", "01111111001100111011", "01001010001100011100", "11000011001101010111", "00111110000100111100", "01001110101100010111", "11000010000101101001", "11010011000100111001", "11011010011011111010", "10110001110100101010", "01010010101101111001", "01000001110100100101", "11000110010101001101", "01100001110100001010", "01010110000101001000", "00110110000100001001", "01001001100101011001", "01001010011100010111", "01000010010100101000", "01000010001101011000", "11001010101100001001", "10111010010111101001", "01000110110100101001", "11010110011100011000", "11000010110100111001", "01000111001100001101", "01000010011100111001", "11001110010100101010", "00110010010100001001", "11000101111100001001",
		 "01001010101100111000", "11001110001100011001", "11000010010100100110", "01001110011100001000", "01001001111101010110", "01000110011100101000", "11001110100101011000", "01001010011100100110", "11000010010101011000", "11001001110110001000", "10111010011110010111", "01001110101100011000", "11010010001100100100", "11000010111100101001", "11011111011100101000", "10111010010100111010", "11100010111100101000", "10111010000100000101", "00111010001100011000", "00111010001100011010", "01000110010100101000", "10111010010100101100", "11000110110100000111", "01000111010100001100", "01001110000100000110", "01000110101100111010", "01010010100100101010", "11001010011100010111", "01001110000101001010", "11000110111100111001", "11001110011011100111", "11001110000100001100", "11001010100101100111", "01001010101100001011", "11000010000101111110", "01000010010101001000", "11011110010100110110", "11000010010100110111", "01100001110100110111", "01000110011100001001", "01001111010100001000", "00111110110111111000", "01010101110100001011", "01001010010101101001", "01001010010100101000", "01000010110100011001", "10111001111100101010", "10111010001101001000", "10110110100100000111", "01000010111100101001",
		 "11001110100100011011", "01000010011100011011", "01010010001101010111", "01000010101101000111", "11000110111100111001", "01100010010100001000", "00111010000100100110", "01001010110100100111", "01110110001110011000", "01000010111100110111", "11001110110101010110", "01001010111100001001", "01010010100100001101", "01001110001100111010", "11010010011101001010", "01001010011100011010", "11000111000100100111", "00111010000101111001", "10101010111110101001", "00101111011100001000", "01001110011110001001", "01000010000100001010", "01000110000110000111", "01000010101100110111", "11011001111100110110", "11010101111100101000", "10110110100100001001", "11000011111100000111", "01010110101110011010", "00111101111100001010", "01001001110101011000", "11000010110101001001", "01001010000101001001", "01000110010100011000", "11000010100100111100", "00111110010100001010", "00111110101100101000", "11001110010110110101", "11101010000101011000", "00111110001011101010", "11001110001100011001", "11011010000100110110", "00111110101101111001", "01010010101101010110", "01011110011100011011", "10111010010110001000", "01100101110101001010", "11010110010101110111", "11010011001101111001", "11001010000101101001",
		 "01000011011101011001", "01001111010011111101", "10111110011110101011", "11000010001100000110", "01000110000100111010", "11000101111100100111", "01000011001100111001", "10111010110101111001", "00111011001100011011", "11001010010011100111", "01011010001100011000", "01111110010101101001", "01011110000101001001", "01010110001101111001", "11101011001100001111", "01100110010100111000", "01010010000111010111", "00111010001100000111", "10111011001100110111", "00110110111100100111", "11000110011100010111", "11010110101011111010", "00111001110110001100", "11001110000101001010", "01000110011101011010", "11001010010100111011", "01010110001101000111", "11000110000101000111", "11011110001011111000", "10111110000111101001", "01001010101100100111", "11010010001100011010", "01001110011100011010", "01000011011100110111", "01011010100101011010", "01010110001100001010", "11001010010101101011", "11001001110100110111", "10111110010110001000", "01000110010100101001", "11010010011100110111", "01000110011101010110", "01000110000100001001", "01001110010111101001", "01001110010101000111", "01000111010100010111", "01001110000101110111", "11000110000110111000", "00111110111101011000", "01001101110110101000",
		 "00111010101100111010", "00111010101100111001", "10111010011100101010", "01000010000101000111", "00111010011101010111", "11001110100101111011", "01001010110101001001", "11010010100110001000", "11000010110100001010", "01010111000100000111", "10110001110100011010", "11010010011110010111", "01011110000100001000", "11000111010100101100", "00111010010100000111", "11100010000100010110", "11000110110100011010", "11001010010101100110", "01011010001100001000", "10111110001100011010", "11001011011100000111", "11001110001100001011", "11000110010100000110", "11001101101100001001", "01010110001110111001", "10111110111101011011", "11001110011110111011", "11001110001101001010", "01011010011100001000", "01000111001110010111", "11001010010100001000", "01001110100100001010", "11000110100100011011", "10110101111100011000", "01000010011100101011", "10111010010100100111", "01111010000101011000", "01001010001111011000", "01000110101100001000", "01000010010100011100", "01001010010100111011", "01001110111100111011", "11100110010100111010", "01000010000101001000", "01010011110011100111", "01111110001101101101", "01100110001100000111", "10111011011011101100", "11100110000100010111", "00110001110101011000",
		 "11001110111100100111", "01000110111101001001", "01011011000101010111", "01011010010100110110", "11000010010100101000", "11000001110101100111", "00111010101100101001", "11001010000101011010", "01000101111110101001", "01000011001101111010", "01000001111101001001", "01010010010100111001", "01010011001100011010", "01000110011100100111", "00110110100100111010", "01010010111101010111", "00110110010100101001", "01000010010011110111", "01001110010101111100", "01001101111100110110", "11100110000100100111", "11101110010100111000", "00111110011101010110", "11010010011110001001", "01001110000100010111", "01001110000100101000", "11001110101100010111", "01001110010110001000", "11000101110011100110", "11000110001100110110", "11011110000101100111", "01001110010100101000", "01001010010100100101", "00111101110100001000", "11000110011100101001", "01000010001101000111", "01001110011100001011", "00110111000011100111", "11000010011101100111", "10110010011101101001", "11001010101011100111", "10111110000100111010", "11100001111110001011", "01001010110100010111", "11001110101101000110", "00111110001011110110", "01000110010101001000", "11010010011100001010", "01001110011100011000", "11000110001100111000",
		 "11001011011101011001", "11000101110111111010", "11000110111011101000", "11001110010100111010", "01100110001011100111", "10111110110100001000", "01011010010100001000", "01010110011100111000", "01100110001100011010", "11000110100101001011", "10111110010100101000", "11010110101101010111", "01001110000100111000", "01111110110100111010", "00111010110100101000", "01011001111100001001", "11010010011101001001", "01101010101100100111", "00111101110100101010", "01001010011100001001", "11001110101100000111", "01010111001100101010", "10111110001100111010", "01000010100100001000", "11000101110101011000", "11000010010100000101", "01000010001100101001", "01000110010100111001", "01011010000100010110", "11000010100110000111", "00111110011100101001", "10111011011100111000", "01001110101101101001", "00111110010100101010", "01001010011101001100", "01010010010100111001", "00111110010100010111", "11000010011100001110", "01000010010100110101", "11100011001011101001", "00111001111100110111", "00111010101100010111", "00110001110100001011", "11001011100011100111", "11000010011100000111", "00111010010100011001", "11010110000100001000", "01001110010101001000", "11001010011100111010", "00110010100101011001", 
		 "11001110001101101000", "01011010101101001000", "10101101100100111000", "00110010101100011000", "00111010011110111011", "10110110001011101000", "01000110110100110101", "10111001111101011000", "00110010001101000110", "11000101101100101000", "10111010001100100111", "01110001111100110101", "11000011111100000101", "11000010011101000111", "00111011001011110110", "01001110010100100111", "01011010101101010110", "00111010000100000111", "00111010011100010101", "00110010000011110110", "11010110111011011100", "10111110011100110111", "01000001110011100110", "00111010001011000111", "01101110010011000110", "11001010000100000111", "10111101110011110101", "00111001100100110110", "01000001110011110100", "10110110000100001000", "11010110000100010111", "00110010000011000110", "10110101011100110110", "11001001100011110110", "10110110000100110111", "11000110010100010111", "01000110010100011000", "11001110011011100110", "00101010001011000110", "00110010000011000110", "00110001111100000111", "01000101110100101000", "00101101111011100101", "11000010010100101001", "11011011100100110110", "01000001111100001010", "00101001110101000101", "01000110000100110111", "00110001110100000111", "11000110011100000110",
		 "01000010011100011000", "10110010110101011010", "00101101101011100110", "11101110101011000110", "00111001110100010111", "01001110000011010101", "00110010001100001011", "10111011001011110111", "00111111011011011000", "11010001101101100111", "01000010000100010110", "11000010000100111001", "00101001011101000111", "10101101111100111000", "01111110000100110110", "11000010100100111000", "00101001000011000110", "01001001100101111011", "11001110101101111000", "10111011000101010111", "01001010110100110101", "01001010010011110111", "01001101100011010110", "10111101111101100110", "00111001110100011001", "01010011001011000111", "01000010011011111000", "10111010101100110111", "10111101110100010111", "00111110001011101000", "11001110011100000111", "10111110010100001001", "10110101100110100110", "11000010000011110101", "01000110011011111010", "11000010100101000111", "00111010010100000101", "01000110010011101000", "11001111001100110111", "11001010000100101001", "01000110011100011000", "01111110000100000101", "10111101011100100100", "11010111001100110101", "01000010010101010111", "00111001111011000110", "01000110010100111010", "00110110000101100111", "01000010000100010110", "11000110000100010110",
		 "00111001110011100101", "00101110000011010110", "01010001110100101010", "01000010000100101000", "10101010000010101000", "01011101111100011000", "01100001101100010110", "00100110110100010110", "00101111000100111000", "00110001110100000101", "11000010110100010100", "11100001110100010101", "01101110101100111001", "01000001111010100111", "10110101110100011000", "00101001111011001001", "01011001111011011010", "10110001100011101010", "10111110010011001000", "00111001101100001010", "01000110010011111010", "11001110101100010101", "01001010101111001000", "10111110011100000111", "01000010010011111001", "00110101111100110111", "00101110001011000110", "00110010011011110111", "01000010000100010110", "00111101011011001001", "01001010010011111000", "01001101110011011001", "00110010001100010111", "01001110100110010111", "10110101110100011100", "10110010010011101000", "10101110100100001000", "00101001101011100110", "10110110111100101001", "11001110001100001000", "01010101100100000100", "01001101101100010110", "00110001110100000110", "10111010011011000101", "01000010001011111000", "11000010011011110110", "01001110101011010101", "11000101111100100101", "01000110110101110101", "10111010010010100100",
		 "01000110011011111000", "00101101110011100110", "10111001100011000111", "10101010101100000110", "11000011110100110101", "11001110100101001000", "11000110010100111000", "11000010010100001000", "00111110001011000111", "11101010010011010101", "00110010001100100101", "01000001110011110111", "00111101101100100111", "11001010010101001000", "01001101101100000111", "10111010011101001010", "10111001100110001001", "11001010011100011011", "01000101111011001000", "11000110000100011000", "01100010000100110101", "01010110100011101000", "01001001101011110111", "10111110101011001001", "01001010100101001001", "10101110011011100101", "10110110010100011001", "11001101100100111000", "00111110110011000110", "10111011001100010110", "11001010011100010111", "10111101100011111001", "11000010011100011010", "00111101111100000111", "01000001111100101010", "10111001111011100111", "00110010010100000110", "00111010000100011000", "00110010010011100110", "10111010100101011000", "00111110100101011001", "00111011000101100110", "10110010011100111001", "10101110011100000110", "11001010000011111001", "00110001111100001000", "01000001110011000111", "11001101111100111001", "10111010000100100101", "00110110011100000110",
		 "10111110001011110111", "00111110010100101000", "10110101110100011001", "00101010011110101000", "01000101010011010110", "11010010011101110110", "00111010110110010111", "00101010011101001001", "10110010101101001010", "11000010100101101000", "11000010000100001011", "00111101111011001010", "10111110001100110101", "11000101101011010110", "10110001101011011001", "01000101100100111000", "00110001110100001000", "01010010010100000110", "01001010111011111010", "11010001111011111000", "11000110100110010110", "00111010001011100110", "10111110010101010111", "11000101010011111010", "00101001111011000101", "10110110010011000111", "10111110010011000111", "11100110011101010110", "00110111100111101000", "01000110110011110110", "10110110110110100110", "11000010011110101100", "10110110000011111010", "10110010011101011010", "00110010110011100111", "01000110011100100110", "10110010100101001001", "10110101111110001000", "10110101100100010111", "01011010110100010101", "00110110001100001000", "11000001110100010111", "01000101111100001001", "00110010101011101000", "10111101110110111001", "01001010011101011010", "00110101110011100101", "00111101110101000110", "00110001111100010110", "10111010011011011000",
		 "10110110010100001010", "10111110001011000110", "00111101111100111010", "10111001011101000111", "00101001110011100101", "10111101111100001001", "00111010000100011001", "10110111100011111010", "00110101111100001000", "10111101010010100110", "00110001100100011000", "01011110011101110101", "11001101111101001010", "10110001100100001001", "10110101100110010110", "10111110010100101001", "10110010111101010111", "10110101100100110100", "10110101111101010110", "11110001100011110111", "10111110100100010111", "10111010011100010110", "01001010001011110111", "11010101100011000110", "10111110010100010101", "10110110010101100110", "11000110110100011000", "00111101111100011000", "00110110011110000101", "11001110011011110110", "01000010101101110111", "10111110000100110110", "01001110010100111000", "11000101110100111001", "10110001111100100110", "00111010001100010110", "01000110011100010110", "10111010000101000110", "11100001111100110111", "01001010010100010110", "10111101111100011000", "11000110011100001010", "01111101110101001010", "01000010011100010101", "01000001110011100110", "11001010011011010101", "10110101101011101010", "01010111010011000101", "00110010011100100110", "01010010101101001000",
		 "01111010000100101000", "01011110011100110111", "01000010101100101001", "01000101110100000101", "01001010001011101001", "01010001111110000111", "01000110000100000101", "10111010110011101010", "11001101101101011000", "10111101101011101010", "10101101111101011000", "10110010100011001000", "10110101100101000110", "00111001111100100111", "10110010011100100110", "01011110001011110111", "11000110000100010110", "01000001100011110101", "11000110000100101000", "00110001101100100111", "01001001101100111000", "00111010011011001000", "01111101110011001000", "01001011000101010101"); 
		weight_ROM(11) <= (
		 "11000001110101011000", "00111001101100000110", "00101001010011001001", "00111001111100000111", "11001011110100100111", "01000110001011101000", "00111001110100100110", "00101101110100000111", "10110110000011001001", "11001001110100101101", "10100110111100011000", "11001010100100111001", "11000010001100000110", "00110010101101010110", "11010010110100111000", "01010010000100101000", "10101110101011100111", "10101010000100000100", "11010110000100000101", "01000011010101010011", "11000010011100010110", "00100010011100100101", "01000110011100111010", "10111001111100100101", "11001001100011110100", "10111110101110010101", "11010010010101110111", "01000011001100111010", "00111101111100010100", "01010010111100111001", "11010010001101000110", "01000110100011000101", "00110010000100001000", "11010110111100000110", "10111110100100111001", "00100101100011101010", "00101101111100101000", "01010110001101100111", "10110001111100100011", "01000010000011100111", "00011001110100101001", "01000110001100010111", "10110101101101000110", "10111010010011101000", "01010010000100011000", "00111110000100000101", "01000110010011111001", "01010101110100000110", "00101010000100010111", "10111010010100101000",
		 "11100011010011110111", "01001001011011101001", "00110001011100000100", "11000001111100100100", "01001111000100110111", "10110010000100000101", "11000011010100110100", "10111001111101000101", "10100110001101101011", "11001011000011111001", "00110010100111010110", "11000110000111011000", "01001001011101010101", "10110010101100101011", "01000010100011110110", "01000010100111010111", "10010110001100001000", "00110010001101110011", "11000101011100111000", "10110110001011011000", "00110010000101011000", "00101010010011000100", "01000010000100101001", "01001010010101001010", "11010011110101010111", "01001010010100110110", "01001010000100110110", "01000110010100111010", "01001001110011100111", "01001001111100010111", "00110101110100001000", "11000011111101001000", "00101101111011101100", "11010010001100110101", "00111110011011100100", "00111001100011111010", "10110010110100000110", "01000010001100000101", "11000010110100110101", "01010110000100111000", "10110001010011111000", "00111110100100011010", "11000010100100110101", "11010110001100110110", "11000010011111010111", "11000001110011000110", "00110010110100000110", "01001110010011100011", "01000110011101011000", "00111010000011100100",
		 "00110010101011110111", "01111101110101011000", "11000010111100100111", "11000011001101110101", "10111001110010111011", "10111010111011110110", "00111001111101101000", "11000010011100011000", "11010010000011110101", "00111010000011000101", "00111111000100010101", "00111010011100011010", "11001110111100110111", "10111111101011111010", "00111110000100111000", "01001110000111010111", "11000010001011001101", "11011010011100111001", "10100010000101001000", "10101110000100101010", "10111110000011010110", "10111110010101010100", "10110110100100010111", "10111010001100011000", "01000111001100010011", "00111010000100100100", "10110010011100101001", "11011001110101000111", "00100010010101000111", "00110101011100111001", "10111010000100010101", "11100010000011110101", "01100110001100111010", "00110010010011110101", "00101101010011000101", "10101110010101000110", "10100101011101001000", "00101010001011110110", "10111001110100000111", "00110110000100110111", "11000010001100010101", "00101001101100000100", "10111010011011100110", "11001011000100101000", "01011110110100110101", "10101010010110100101", "00110001101011000100", "11110010000101110100", "10110010010011110110", "00101101101100110101",
		 "00111110000100101000", "10101101101100101001", "11000010010101101001", "10100010000100110101", "10111010010011100101", "10111110101011110110", "01000010011100011001", "00110010000100100110", "01010010000101011000", "10110001110100000110", "00110110001100000110", "10111010011100000110", "00101101111101100100", "11000010001011100111", "00110010101011110101", "10111010010100011100", "11000010111100011001", "10111110000011110111", "01000110011101010111", "01000110011100011010", "11000110011101110101", "10101110010100001010", "11000110110100110111", "11001110111011100110", "10110110000111110111", "10101101111101111001", "00100001100010100111", "10111010010100010111", "00100110010010110111", "01000001101101000111", "11001010001110010100", "01001101110011101001", "00111001111101000111", "01000001111011110100", "10111010000100110110", "10111110101101000110", "01001110101110111000", "01010010110011100100", "10110010001101010101", "01001001111100110101", "00111010110100010110", "01000010011011100110", "10110101101011110110", "11100010110100011010", "11011110010011110101", "10110001111100101000", "10111110010010100100", "10101001110100101000", "00111110100011000110", "10110010001011010101",
		 "01001110000100111000", "01001010100100000100", "01001001111100111100", "01001010010101100110", "01010011111101110101", "10101001110100100110", "01010010001100011000", "00110110011100001000", "10110110100011100111", "01000001101100111000", "10111001101100101000", "00111101111100000110", "01010110001100110110", "11000110011011101000", "10110110001100100111", "11001001110101010101", "10110001110100100111", "11001110010110110110", "11011010010100110110", "01010010000110101001", "10111110011100010111", "01100110101100111000", "00111110100100110011", "10100001100100101000", "01001010011101110111", "10100101111100010101", "11100001111100011001", "00111001100111010111", "11000110001101001001", "01001010011100010111", "10110110010011010111", "01100110000101111010", "10111110001100101001", "11100001111101101001", "00110010010100110111", "10110010101100100110", "00111010000011001001", "10110110010100111000", "10111010100100111101", "11101010000100100111", "00111001110100100100", "01000010001100010101", "00110101111100000111", "10111010001011010101", "11000011001100110111", "00111010000100000101", "11001101110100010110", "10111110010110111011", "00111010001100000101", "01000110000100111000",
		 "01101011000100111011", "00111101100101000111", "11001101011101001000", "11000110000100100110", "00101001101100101000", "00110001101100100111", "10111101110100001010", "00111011011011100111", "00100101110101010101", "11000101110010110110", "10111010101100011001", "10111010011011011011", "00101101110101101000", "11010010010100001000", "10101101110100010101", "00101111100011111011", "10110110001011111000", "10110110001101000101", "01001010010111111010", "00110010000101010101", "00111010111101010111", "10101110100101001011", "00110101110011010111", "01010110010011010101", "11001110010101010110", "11001010000100001001", "00101001110100001000", "00101001100100110110", "11001010010101010100", "01000110011011100100", "10111110011100010111", "01000010001100110100", "11010001111011110101", "01001111000100100111", "00101010000011000110", "00111010101011110110", "01001010010011110111", "01000001110011110101", "01111110100100010110", "10110010000101000100", "10111101111100010111", "10110010011101011011", "00110010110100101001", "01001010010111010110", "00111110010101100110", "01000110000101100101", "10110010010100001001", "00110111001011100110", "01001111011100101010", "00011001111110011000",
		 "00111101110100010101", "01000010010110011000", "10101110000100110111", "10110101010100010100", "11001010001100111010", "10110110101011101000", "11001111010011110110", "00110010011100101000", "01100101101100101000", "00111001111011101010", "10100110011100100111", "10111010110111101111", "01001010011101010111", "10101010100101100110", "11010110111100110111", "10101110001011100101", "00101001110100100110", "10101010001100000101", "10111110011100101000", "10101010111011101000", "11001011010100101000", "00101110011100000101", "00100001110011111001", "11000001101100000101", "11000010100011110110", "01000001111100010100", "10111010001100001000", "10111110100100000110", "00101101010101010011", "11010110010100111000", "10110001100100100111", "00111010011110010111", "00101010100100000101", "11000101110011111001", "01000110010101110110", "01000110000011110110", "10110001110100010100", "11001010001100011000", "01001011000100100110", "00110010101010110110", "00110010001100100101", "11101010011011100110", "10111110110011100111", "00110010010101010111", "01001110100100000110", "10111010000100011000", "11001001110011100101", "01010110000100010111", "10110110010100111001", "00111101110100010101", 
		 "01100010000100011001", "11000101111100101001", "10110001111011111000", "11010010001100111000", "01111101110100000111", "10111010110100000111", "11000010010011110011", "10110110000011101010", "10111001111100010110", "10110010010101111001", "00110001110011101001", "01011010100100100110", "10111010000101010110", "00110010011101101000", "11010010100100011010", "01001010010100100101", "00111110010100001000", "01000110010101111001", "01010110001011110101", "01010110010100010111", "01101001110100111000", "11000010111100101000", "01000110011100010110", "01001010001101000011", "11000101011101000101", "01100010010101010110", "01000010101101010111", "10111110001100111010", "01111010010100100110", "00111001101100101010", "11001110111011111101", "01001111001010100111", "10111010010100100101", "00111010011101110101", "00111010110100101001", "10111111010100010110", "01001010010100110111", "00110110110110000101", "01000110010100100100", "01001001110101001001", "01001110001101001001", "10111101111101000111", "10110110001101001000", "01000110011100001010", "11000101110100101001", "10111010010101110101", "11011010000100010111", "01001110011100110111", "00111011000101001001", "11000110000100011010",
		 "11001110001011111000", "11001011001101101000", "00111010101110101011", "00110010011011001000", "10111110011100011001", "11001110001101000111", "11000001110011010101", "11011001101100000101", "00111010001101111000", "10111010010100010110", "11000010011100101000", "01110110011100010111", "01001110100100010100", "01001110010110100110", "00111010000100111001", "11010010000100010111", "10101010101100001010", "01000010101101011010", "00111010001101011100", "01001010001100110111", "01011010101100111000", "11101010001110010100", "11001010010101111000", "11001010000011101000", "10101010001100010111", "01000110011100101010", "01000110010011010110", "01011010000100001101", "01011010000100011010", "11001110011101010111", "11000110100100111010", "10111101110101111010", "10101110001100001010", "01010110110100011000", "01000010001011100101", "11100110001011100111", "11001010001100010111", "11000010101100000110", "11010110100100110111", "10111110100100001000", "11100001101101010110", "01001110010101000101", "11000110011011101011", "01111001111100111000", "10111010100100101000", "10101110011011001001", "00111010001100001111", "11001110000100010110", "11000110101100001000", "00110001110100010111",
		 "10111010101101100111", "01001110101101000110", "00111011011011001001", "01110010000100100101", "11001010101100111000", "00111010011011100100", "00110010110100011011", "00100010000100100011", "01000101111100010101", "10111110000011110100", "01000110000100100101", "01000110001100011000", "01010110101101011000", "10111010101101111000", "01000001110101101011", "00111110000100100110", "01001010011100100111", "01001010000100001000", "11000010010011100111", "00111010001100111011", "11001010100100101000", "11001010110100110101", "10110010001110101000", "01000010111011101001", "10111110110100100101", "11100010101100100111", "11000001010100001000", "01001101011011110100", "11010110011100000111", "10011101111100001010", "00111101110101010110", "10111110010101010101", "01001010000100000111", "10110110000011110110", "00110010000100001000", "10111101100011101011", "10101001111011100111", "01010010000011110100", "01101010010101011000", "01000110100100101010", "01100010011100000100", "11010011001011110110", "00111010100100100110", "00110111011100001000", "11001110000101010111", "01000001111100000100", "00111110000011101000", "01011001110100010111", "01000001110011100110", "10111110010100010110",
		 "01010010011100001001", "10111110100011100101", "10111101111101001000", "00100010011011100101", "01100011011100000110", "11000110101100000110", "01000111010100110111", "10110110100011101000", "11100011001100110111", "00110010000100001000", "00111110101100110110", "11001101111101100101", "10110101101101100110", "10110011100100101000", "11010110001100010011", "10111110010110001001", "10110010100100011000", "11001101111100111000", "00111001111100010110", "00111010100100010110", "10111110110101010110", "00111001110110011000", "11010010100101000111", "11010010011100001010", "10111010110011111001", "10100101110101011001", "00101110011011101001", "01010010010101010110", "10110010010011001011", "10110110010100100111", "01000110111100000101", "11001110000100011000", "11011110001100000111", "01000010101011110110", "00110010001011100100", "00111001101100101100", "00111010010100111000", "10101110010100101111", "01001110000011100101", "01001010010101111000", "00110001110011110100", "00111110000100010100", "10111110001110011000", "11000110010100110101", "01010001110011101000", "01001010000100110100", "11000010010011100111", "00110111100011111001", "10111110111100101110", "11010011011100000111",
		 "01010110010101011000", "01001010000101000111", "11001010100100111110", "00111010010100111000", "00101110100100011000", "10110001110100000111", "01001010010100010111", "00110110001101000111", "10100010110011011001", "11010110111101001001", "10101010000100011011", "10110010011100111001", "11000101110101011011", "11000010001100011010", "00110010000100011010", "10111110001100010110", "01000010111100011011", "00111010001100010011", "00111010111100010101", "11000111001101011000", "10111110011100001001", "11000011011110011010", "11001010001100010101", "00100101100100110111", "10111010010011010101", "10110110011011110110", "00110110011100001011", "10111001111100001000", "01001110010110001001", "11001010111011100111", "00101110100101011011", "01000110011100111001", "01101110011100111001", "10111111000101101000", "01001010010100110100", "11000110010100010101", "10110001111010101100", "11000001111100101000", "10110110001100111000", "00111010000100010101", "10110110011100010101", "01001011110100111010", "00101001101101110101", "01001111011100001001", "11000110000100101111", "11010011011100000111", "10101101110100100101", "00111010100100011010", "01001010011011010111", "00110010000100111001",
		 "10111010010100010111", "00111001110101001011", "11001010010011101000", "11010110101101011000", "00110001100100111000", "10110010100100111000", "11100010001100101000", "11001010001100111000", "00100111000011101000", "10111110010011101000", "01000001110100100111", "10111010001100001000", "00111110111101001001", "11001001101101001110", "10110010000011110100", "11001010001100111010", "00101011011100101010", "00110001110011101001", "11000010101011110111", "01100010000101001011", "10111010001101011000", "10111001111100000110", "01001101111011100111", "00110101110011100101", "00111110110011101111", "11000011000100100111", "10111101111100001001", "10101101110110111001", "00111110001100000111", "11000110100101000101", "11000010101110111001", "00111010011100000101", "11011110011100100111", "10110010101100110111", "10110010001100100111", "11000010010100011001", "01010110110100101001", "11001110001100000100", "00110010101011100101", "10100110100100001011", "10111010000100001011", "01010111010011101000", "00110110010100100110", "00101111101100000111", "10101010101101000100", "00111010010011100100", "01011011001100101000", "00101001110100000101", "11000010000101101010", "11001111000100000111",
		 "11110010001100100110", "01010110001100111001", "00111110100100011001", "10110101110100100111", "11001011011100010101", "00101010010101111010", "00111110111011010110", "11000110011101100111", "10111110011100001000", "10101010000100011001", "00101110001100100111", "01001011011011001001", "11100110001100000111", "10101010100100001000", "11001010010011111001", "00110010110111110011", "10111101111100011001", "10111110010100010111", "00111110100101001010", "11000010000110001000", "11000010000100101000", "00101010000101100111", "00111101111110001000", "00110010000100101000", "11000010000100000110", "01010010111101010101", "00110110010011110101", "01000110001011110101", "00111001100100010101", "00111110000011111100", "11001110011010100111", "01100101110100111001", "11000110101101000101", "11000110001101110110", "11000001110100110111", "01000110000100100111", "11010010100100110110", "11000110100011101001", "00111010010100010101", "10100010010110001001", "00110010011011111001", "00110010100100110100", "00110010001100100110", "11011110001100101010", "01001110110101110101", "11001110101101001001", "00100010001100010111", "10111010011100111010", "00111010001011100100", "00100001101011000101", 
		 "10111010101101001010", "11000101010100001000", "10101010001011010111", "10111110011100111000", "10100110000100011010", "10101101011100001000", "00110110000101000110", "00101110001100001100", "11000110100100000101", "10111010100100111000", "10100110000100001010", "11101110000011000110", "00100001011011100100", "01000010011011100101", "11010110100101000100", "01001110001100001001", "00111010011011110101", "00101110101101110101", "01000010000101010101", "00110110010011110100", "00111110011011110110", "10100001101011101001", "11001110011100010101", "10111110011100111110", "11001101110100000100", "00111010000100000110", "01001110000011110101", "10110001110101000111", "10110001111101010011", "10110010011100111000", "11101010110011110110", "01000010001010110100", "00110001110011100110", "00101110010100010110", "10101101110100110111", "10011010011100001001", "00110110000100110110", "10110111010011000011", "10100001111100000100", "00111010011100100011", "10100010010011100110", "11000010000101000101", "10100001100110100110", "10100001111101000110", "01000010011101011000", "00111110100100010101", "01000010001011100011", "01100110100110000110", "00100001111100000110", "10101010010100101000",
		 "11000101100110101010", "10101101110100111001", "00111101101100111001", "10101010110011100101", "01000110000100000101", "01000010000100100100", "10111010000100010101", "01100010101110010101", "00110010000101000100", "10110010011100111000", "01001001110101110100", "00111110000101000110", "01000010010011010101", "11001001100101011001", "01000010000100010110", "11001010101100110100", "10110101110011100110", "01001010111101010100", "10101101101110000110", "10111010010011010110", "01010010011100101100", "01001010010100010111", "11001010000100000110", "10101010000011111000", "10100101110100010101", "11010110000101010111", "00111010000010110101", "01001110000110010110", "01010001110101000111", "11100110000100100111", "00100010101100101000", "11000111001101010110", "00101101110010111010", "01100110001100001010", "10110110010100000100", "00100010001010100101", "10101101100100100010", "00100010100100100101", "01000010010100010101", "01000010000011101001", "10110010110100110101", "10100110010101000110", "10110101101100010111", "01001110010100010100", "01000010000011101000", "10111011010011100100", "00110010100110100101", "10101010011011100101", "10111010010100101001", "00110010000100000101",
		 "10110001111011110101", "00110001111100100100", "10101001100100100110", "10111010010011101000", "00111001100100001001", "01010010001011101000", "00111110000100100110", "10110010000101000101", "01000110000100100110", "11000010000011100111", "00110110100100010101", "01001010010100010110", "11010010011100001010", "10111110011011010111", "11001110010100010110", "00111010100100100101", "00111011001011110101", "10111010010101101001", "10100010001011110110", "10101101010100000111", "00110101110110001000", "00111010001100000100", "01000010011101001000", "00111110000101011000", "10111010010011100101", "11000010001101110100", "11001101110101100111", "11001001101011110110", "10101110000110100101", "00011101111101011000", "01000010100101110101", "11001010000100101001", "11100110000101010111", "01010010000011010100", "01001101101110000110", "00100001111100110101", "10110110000011000111", "01000110100011100111", "10110001111100101001", "10111010010111100101", "10100001101011100011", "00110001011100000100", "10110001110011100100", "10110001111100000111", "11001110100100011011", "01011110101100010101", "00101101100010000110", "00110010101100101000", "01010110010010110101", "10110101101100100100",
		 "01010010011010100111", "00110001011100100110", "10101110011100101000", "00110011110100000111", "11001010000110011001", "00110001100011100101", "01000110101100010111", "00100010010011100101", "11000110001100010110", "00110010010011100100", "00110101100100010011", "11000110000011100110", "00110001100100110100", "11000110000011110111", "00110110001100010011", "11000010100011011000", "10101110110100000111", "00111110000100000110", "00100010000100000110", "10100101101100101010", "00110001111100110100", "11000101110011101000", "01000010011100001001", "01010011001011111101", "10111010111011111000", "00100010010101001000", "01101101100010011000", "01001010100011110110", "00111110100011010101", "00100011001011111000", "10110001110011100110", "01100101100011010111", "01010010001100100111", "00110010001100111001", "00101110000100000011", "00111010001100110110", "01001101110100111010", "10101010000011100110", "10100101010011110100", "11010110101100010100", "00101001110011101000", "00111110001100000101", "11001101011100001001", "11100010011011100110", "00110101011011000101", "10101001111100010101", "10111001110010100100", "01010001110100101000", "10100101111101001000", "01001011001010100101",
		 "11001010011100111011", "01000110101100000101", "01000010001101011010", "01001101111011100100", "10111110100011110011", "10111010000101100100", "01000110001100110101", "00110110000111110111", "10110110101100010110", "00111001101011000111", "00011001100100000111", "00110101110010110110", "10111010010100110101", "01011010100100100111", "10110010000100000111", "01000101110011110111", "00101010000011100111", "00101001110011110100", "00111001111011010111", "01000010101110101001", "00110010011100110111", "10101010010101000101", "00111001100011100111", "11000110000100001000", "00101001011011110101", "10101001111011100100", "00101101010100111001", "10110101001100110101", "01011110000100110110", "00111110011100111000", "00110110000011000111", "01001110010100010111", "10111101110101111000", "10101110011100101111", "00011110101100010110", "10111001111010110100", "10101001100011111101", "00100010001100000110", "10111001101100010111", "00110010000011100101", "10111110011101100110", "11100010010100010101", "11001001101101001000", "10111010011011110110", "11000110001100011000", "10110001111011000110", "00111001010100010111", "10111010101101000111", "10110001011100100110", "00101010101100101010",
		 "00110010100101011001", "10100101100100110111", "01000110000101101001", "00101010101100100110", "00110001010101000110", "10111010011100000111", "01011101111101110110", "01001011001100001001", "10101101100100010101", "00110101000010111011", "01010110111101011000", "10110110011100110101", "11001010001101011011", "10101010001101101000", "00111101111100010111", "00110110010100101100", "00101010011011110101", "10100010001100011010", "10110110001101010110", "01010010100100110011", "01000110100101010101", "00111010101011110110", "10111001111100000100", "11000001010011011001", "00111010010110010101", "00101001110100001000", "10110110001100101001", "01001001101101100110", "11001001101100010101", "00101110010100000100", "11001010010100110110", "10011010001100010011", "10110010101100111011", "10110101111011111000", "10110010100101111001", "01010110010100000111", "11001010010101010111", "00101110000011110110", "11000010011011110101", "10110010000100000101", "10110101101110010111", "01001010011011100111", "01000011000100000111", "00101001111011110110", "10101010011100010101", "10100010011100000010", "11001101111011011001", "00100110010100100101", "01011010011100011001", "10110001111101011100",
		 "10111011000100010101", "00110001110100111010", "00111110111100010110", "01001001100011000011", "00111001100011110100", "10100001111100000111", "01000101011011110101", "10111101111100011001", "11000101011100010111", "10101101110011001001", "00110010010100110110", "00110101111100111000", "10110011001011110111", "10101001111011100100", "00110101110101100111", "01000010101011111000", "11001010000011101100", "10101010000100010101", "10111101111011000111", "00101001100011010101", "11010110000011111000", "10110010111011000110", "00110010010100010110", "01000001000100110101"); 
		weight_ROM(12) <= (
		 "10111101111101101011", "11100010011110001000", "01000010100100001001", "01000010001011101000", "01000110100111001000", "10110101111101001000", "11001110110100010110", "11011010010101101000", "00100010001101100110", "11000010000101011000", "01000010010100001000", "11000110001100010110", "01101110011100101001", "11010110100100011000", "00111110001100010111", "11000110100100101100", "00110010111011101000", "11010010101100110111", "01000110001100000111", "01100001110110110110", "11001010001011100101", "10111110101101001001", "11001010000100000111", "00111001111100000110", "11011101110100000110", "11000011000100111001", "11001010010100110101", "00111001100100010110", "01001010010100010111", "10111101100100011001", "01010110001100111000", "00111010010100000111", "10110110000100110111", "01000010001101001001", "11010111100100110111", "01011110000101010111", "01000010000100100111", "01001010011011110111", "01010110010101000100", "00110010000100100101", "00110101111100101000", "00111010000101100111", "00111101101100100111", "01001011111101000110", "11000110000100011001", "11010010000101001000", "00101001111100000111", "00111010000011111000", "00101001110100111010", "10111010011011101000",
		 "01010001111100111001", "10110010100011101011", "01100101111100111000", "01011110111101000111", "01001110110101010110", "00111110000100010110", "01010110101100001000", "00111010001100010111", "11011110100101110111", "11110010001011101000", "11000110010100010111", "01010001111100011000", "00111001101100101101", "10111010010111111000", "01001110001100101010", "11011010010101000111", "00101010000100100111", "01001110001111000111", "00110001110100111001", "11010110010101001110", "11001010000101010110", "00111010100110000110", "01010110100101010110", "10110101101011010111", "00111001110011001001", "01101110011011101010", "01001110100100011010", "10111110101100011000", "11001110000100101001", "11011110101101010110", "11011010010101100110", "01010001111101011001", "10110101101100100110", "11100010000011100110", "11000110011100110111", "01001001110100100111", "00111010100011100111", "01000111001101101000", "11000010111100011000", "11010010101100101010", "01001001111101111000", "11011110100100111101", "11010010011011100110", "01010010011100110110", "01010011000100010111", "11000010011101011011", "11000010000100001111", "11000110011101011010", "00111001101100010111", "10111010000100010110",
		 "01000010000111100110", "00111110000100000101", "01000010100110001001", "00111010000100001001", "10110101110011100111", "11001110010100111010", "01011010111101000110", "00110010100100100111", "01000010011100010101", "00111010110100000101", "01000001110100010111", "11001010001100111000", "01001110011011110111", "00110110000100001001", "10111010011100101111", "01000010101100110110", "01001010001101100111", "10110001110011111010", "10111010011101000111", "00101110001011100111", "11011010100100001000", "11000010000100101010", "01001110001100001000", "10110010010100101001", "00110110110100101001", "01000010011110011001", "00110110001011000110", "00111010010100011011", "11100110001101001000", "11011101101100000111", "00111001111101011001", "01001101111100111001", "00110001111100000111", "00111001110100010111", "11001110000100111011", "10101110010100100111", "10110001100100001010", "00111010011100101000", "11001110100110001011", "11001110010100101001", "01001101110011101000", "00111110101101011000", "00101010010100000111", "01011110001101000110", "11010001111100000111", "01010010110100011001", "00111010011100000111", "11011010011100000111", "11011110110101010101", "00111010000100000110",
		 "01101010011011111000", "00111011110011001010", "10110001110101100111", "10110010101101101101", "11000010100101000110", "11001010011011000111", "01000010011100110111", "10101010000100100111", "11000110100100111001", "11011001110011111001", "01010010011100100111", "00111010000011100110", "00111101101011100110", "10111110000101011011", "11001110001101011001", "10110010100100101001", "10110010101100101001", "11001110101101001001", "01000110010100011011", "11001110101100001010", "01010010010101110110", "11000010001100101001", "01001010001100101000", "11000110100100101000", "11000110000100001110", "01000101111101000111", "10111110000100110111", "11100010100111111010", "11010011001101010110", "10110010000101010111", "01001010000011110110", "01010101110100110110", "01001001101101001011", "01010010001100011001", "01010001111100000110", "01000010001101101000", "11000110100100000111", "11001010000110100111", "00101001010100000110", "10111110101100011000", "01000110000100101001", "00111110010100000111", "11000010101101000111", "10111010000101100111", "00111010000100011000", "01000110101100001001", "00111110000010111001", "10111010001101111010", "11011010001100000101", "00111110000111100111",
		 "11010010101100011001", "01000010000100001000", "11000010101100011001", "00111010101110101010", "00110110000101000111", "11001010001100111000", "01000110000100110111", "11100010000011111001", "10101010100100011010", "01011010001100100111", "10111010100100111000", "11000010100011111000", "11010110010100010100", "01001010001100001010", "11000011000101001001", "01001110011100110111", "00111010001100101001", "01000110011101010111", "11000001111101001001", "01010010011100001001", "11001111001100111001", "01000110111100010111", "01011010001101010101", "10111101111100111011", "00111010001011111010", "10101010010100100110", "11001101110011100111", "11000110000100110111", "11001011001011101000", "01000010001110110110", "10101010111101000110", "10111110010100100111", "10111110000100001000", "10110101110100001010", "01000110000100111001", "00111010100100000101", "10111110000100001000", "10110010111101011000", "11001110000100001010", "01010110010101110111", "01000010001100111001", "11001110000101010110", "00101010001011101000", "00111010110101101010", "10111110011100101001", "11010010000100110111", "11000010101100100110", "11001110001100101100", "01001001111011110110", "10110010101100011011",
		 "11010010001011101001", "01000110001100001001", "00111001111101000111", "01001110011101001000", "00110010000100000110", "11000010100110111001", "01100110101100101001", "11001110100100101000", "01100010000110101000", "11000110010011001010", "00111001110011011110", "00110010101011111000", "11001010101101000110", "01010010000100001011", "11100110010101001000", "01001101110100001001", "11001110100101010111", "11011110001100101011", "10110110100011111000", "01000010000011011010", "11000110001110110101", "11000010001101001000", "00110110000101000110", "00111001100100000110", "11001010011101001001", "11000110010100011100", "11001001110110011001", "10110110101100001000", "00111010011101001001", "11000010001100000101", "01001010010100100111", "01010010101101010111", "11010010010100110111", "11010110000011101000", "10110010001101100110", "00111110001100110110", "01000110111111001111", "01010010101011100111", "11010010111011010110", "11010010000011101001", "10111011111100111000", "11000110100111101001", "10111110010101100111", "01000110001100010111", "01000010100100000111", "11010010011100010110", "11000110001101011010", "01001001110100100111", "01000010011100101000", "01001001111100111010",
		 "11000010001100000110", "10111110101110111000", "01001010111101011001", "00111101100011100111", "00111110001101010110", "00111110011011101000", "11000110100011100111", "11001110100100001000", "10110101010101101001", "10110110001100101100", "10110110000101101001", "10111110010100000110", "01000110101100010111", "10111010111100000111", "00110010111101101000", "11001110001011110110", "11000010001101111000", "00111001110011110111", "00111110011011101000", "11001001111101101010", "01000010001100001001", "00111001111100001001", "01000101110011101000", "01001001111100010111", "11000011001100011000", "01000101110101110111", "11010110101101010101", "01000111100100011000", "11010110111101101000", "01000011010011101010", "11000101101101000111", "01000110000100101011", "10100010101100111000", "01000011000100001001", "01010110010100010111", "01010101110011110111", "11011110000100000110", "10110010111100111000", "01000010010101010111", "10110010011100101000", "00111110010100111000", "01001110010011110110", "11000001111101000111", "11010110101101101000", "01010110100100011000", "01001110101011101001", "11000010010100001000", "10111110001101111001", "00111111001100100110", "00110110010100111011", 
		 "01000011001100101000", "11000011110100010111", "11001110100100110111", "01000110000100001010", "01000110010101011000", "00111110001101000111", "11001110100101011001", "10111010010011111000", "11000001110100101000", "11001110101101001010", "11000010100100010111", "11001010100100100111", "11010010101100100110", "11101010011100001000", "10111010000011110111", "01000010010111110111", "00111110001100111001", "11000001110100111000", "11000101110101011001", "10111010010100110111", "11001011010100001000", "11010110101100101001", "11100110000100000111", "11011110001100111000", "11010010110011110110", "11000011011011101000", "11010110010100111001", "00111110010011101000", "11001010101101111000", "01010011010100001000", "01010110110100101000", "01000110111100101001", "11001110101100100111", "11001110101100101000", "01000010001100001001", "01100110101011111000", "01010010000100011001", "01001010101100101001", "11000011111101011001", "01010110100100101010", "01000110110100001000", "01001111010100001100", "01000011001100011001", "11010110010100101010", "11001010100100001001", "11011010000100010111", "01000111010011101001", "11000110011100011000", "01100110000100011000", "00111010100111011001",
		 "01000010010100100111", "11000110000100001011", "11001010010101011000", "11010001110100111001", "11010110010100001001", "01011010001101010111", "11010101111101110111", "11001010111100111000", "01100010001101001100", "01000010011100011000", "00110010000100011001", "11000110111100111010", "11010001111101000110", "11000001111101111001", "01001010110100101110", "11010110010100011010", "01010110101100101001", "01000110011100111000", "11001001111100100111", "01000010110100101000", "00111010011101111001", "11001110000100001001", "11000010001100001011", "01000110001011101001", "11001110010100001000", "01010010001100001010", "11001010110110001001", "11000110010110001001", "01010110111101011010", "11100010000100101111", "01000110011100011110", "01010111101100001010", "00110110001100001011", "11001010010100111101", "01000001111100001000", "11000110101101001000", "01101110001100111000", "01000110110100101000", "11010110001100101001", "11010110001100001010", "11000010010100000111", "11001010010011101001", "11001110101100011010", "11001010100100111011", "00111010000100101001", "11100010111100111000", "11100010000111111000", "11010010001100111000", "10111010000011101011", "11010010000100000111",
		 "01000101111100001000", "01001110010101110111", "00111011100101001001", "00111010100101001000", "11000010001100101001", "00111110100100000111", "11101110100111101010", "01000110100101011101", "01001110010100111011", "11001110111100110111", "11010010011100111000", "11100110011101001010", "11010110010100011011", "11000010001100011001", "01100010001100011001", "11000010101100001000", "01010110010100110111", "11001110001100100111", "11001010000100111000", "01000101111100111000", "01000010010101011001", "01001010011101001010", "11001110010101011010", "00111010110011111001", "01000010000110001001", "01001110100100100110", "10111101110101101010", "11010001100100001000", "00111110001100001000", "01000110101101111001", "11010110101100010111", "11000101111101001000", "01001010100110011110", "11001010100110011010", "11001110010011111001", "10111110100100101001", "01010110000100011001", "01000110010100101011", "01000010010101000111", "01001010000100110111", "11100110111100101100", "01000010100100111001", "01001110101101011010", "01001011010100111000", "11001010110101111010", "01000010001100011000", "01000110010101100111", "11100010011100001010", "01000001111100101000", "01100010101100111010",
		 "11000010101100111001", "10111010100100101010", "11000001111110011001", "11010110111100011010", "01011010101100111000", "00111011111100011001", "11000110011110010111", "10111110010100111001", "01011110001100111001", "11001110100100100111", "01001110000101001001", "00111001111101111000", "11101111001101101000", "01000111001100011000", "11010110010100111000", "10111110000101111010", "11100001110101001000", "11000010011100100111", "10111110101100101001", "10111110000011101000", "11000010101100111001", "11001110000101011010", "01011010101100011000", "11001001111100001001", "01101010010101111001", "01100101111101001011", "01100010001100001001", "01000101111100110111", "01001001111110000111", "00110010000011111000", "11000011010100111001", "01000110010110001011", "00111110101100111000", "01000110001110111000", "01001010001101011000", "01101110101100011000", "11011001111011111010", "11010010101110011010", "11001011101101111000", "11001110100100101100", "01111011000100111000", "10111010001100011001", "11001101111011101001", "11001010000100101000", "11010110011100111001", "00111010000100000110", "01000111001100101101", "11001111001100011010", "00111110010100001001", "11001010100100111001",
		 "11000010001100111100", "11001010010100001010", "01001110000011111001", "11001011000100101100", "01001010000100011001", "01001101111011100111", "01000110101110111101", "01001110001100011010", "01001110001100101001", "11000010100100011001", "11000010011100001100", "11000111010011101001", "01001110111100001001", "11000110001100001010", "11000010000011111000", "11000110000100000111", "01001111010100101000", "10111110110100100111", "11011010010101111001", "01001010011100101011", "11001011001100011010", "11000110001110101000", "01000010010100101001", "01000110011101101111", "11001010010100111001", "11000110011100111000", "11010110011100101000", "01001110001100101001", "11001110010110001100", "11001110010110011010", "11000110010101011001", "11010010001011101001", "01000110011101101101", "10111010011101001001", "11001001111100001001", "01110011000100001000", "01000001111100011011", "01111110111100000111", "00110111000100000111", "01011110100100111000", "01001110000101100111", "01111110100100111000", "01000010001111001010", "11001110000100111011", "11010010011101001000", "01000011001101011010", "11010001111100101010", "00111010010100011000", "11001010001100111001", "01001011110100011000",
		 "01010010001100101001", "01000110101100111010", "01011110011100001010", "00111010001100101011", "01010110011100101001", "01010110011101101001", "11010110100101101010", "11010110011100101010", "01000010000011100111", "11010001110011111001", "11001110011111011001", "10111110001100011001", "00111110001100011010", "00111110110101011001", "01001010001100111000", "01001110010100111000", "00111010000100111000", "11001010010100000110", "11011110100100101111", "11001110000101010111", "01000010000100011100", "01011110001100000111", "11001010010111101000", "01101010001011110111", "11001010000101001011", "11001010011101011001", "11011110011101011010", "01000110010100111000", "01000011000100011001", "01100010011110101011", "01001110011110101010", "11010010001100111001", "00111110100100101001", "01000110011100011001", "11001110111100011011", "11001110000100011000", "01101010111110011000", "01101010001100000111", "01101110011110010111", "01000110001100001011", "01011001111100111001", "11100110001100011001", "10111010001100111010", "10111110111100101001", "11110110010100111000", "11000010100101011001", "01010110000101011000", "11100110000100011001", "10111110010100001001", "11000001110100011000",
		 "01110101111100101001", "00111001111100111001", "11001101110111001000", "11100001110100111000", "11011010000100111100", "01001010101101001011", "01100010100111101010", "01000010000100111011", "01000110001110011110", "01010010010101001001", "11011010010100000111", "01010110011100111001", "01110010011100101001", "11001110010101001000", "11010001110011111001", "11011010000100101011", "01010010010100111001", "01000110100101101000", "10111110000100011000", "11001010101100101000", "11001010010101010111", "11000101111100010111", "11000110001100111000", "01000110001100101000", "11100010010100101000", "11001010010101010111", "11001110001100111000", "10111010010111101011", "01001110100100111000", "10111010010101101001", "01001110000101011010", "11001110001100101001", "01000101110100101001", "01001110001101011000", "11010010100100011000", "01000110110101011000", "01010110000100001001", "01010110000100101000", "11000001111100001000", "00111110001100011001", "01000001111101101000", "01001110101100111011", "11001010100100101001", "11010111010101000111", "10111110111101001010", "11001001110111010111", "11011111011101011100", "01010101110111111110", "11001010101101011000", "00110110010100111011", 
		 "11000110000011111011", "01001010011011100111", "10110001110100111001", "11000110010111001001", "11000010100100001001", "10111010010101101100", "00111110000100011000", "00111010000100011001", "00110110101100101110", "00110010100011111000", "10101010010100001000", "01000010001011100110", "01001101110101000100", "11010010001100000111", "01000110101101100111", "11000010011100001010", "01011110101100111000", "00111101110100010110", "00111110100101000111", "00111011011100110110", "01111010010100011001", "10101001101011101000", "01011110110100111001", "00101010010101111000", "11000101011101010110", "00111010110110000110", "01010010001110010110", "01010010000100111101", "10111010000101110110", "10101010000101001011", "11001101110110011000", "11011101111101100111", "01000101110100010101", "11001010111100110110", "11000010011101011010", "10110010010100001001", "00110101110100111000", "01000110100100000101", "10110110011011100101", "11010010111100000101", "10110001011110000111", "01000010010100001010", "11010010101100001001", "10111010001110111001", "11101010100100011000", "01010110011100110111", "01000011010100100101", "11000110000100001000", "00111110011100111000", "01000110100100100111",
		 "11101110000100101000", "11001110101101101010", "11001001110110000101", "01011010011011001001", "11001010100100110100", "11010010010110000111", "01001110110101110110", "01001010010101100110", "11101010001101110110", "01000010001100011001", "00111010001101101010", "00111110000101101000", "11001110110101110100", "01101010011100111001", "01000010101100011000", "00111010101100010111", "10110010000101001001", "11000110000100101000", "00101010011100001010", "01010110010100011001", "01010110101100110111", "01001101111100110111", "01001010001101001000", "11001001101101001000", "00110110011100000100", "11100110000100101001", "11000010011110010110", "01001110010100001000", "11000110011100010111", "11011010100100110111", "01000110000011111000", "11001110011101011000", "00100110000100100111", "11001010101100101011", "01000110000100001100", "01000110010101100111", "10110101110100000101", "11011111011011100110", "10111110100100011010", "10111010011100111000", "10111110000100010111", "01001101111100000100", "01001101111100101000", "11000110001101010110", "11000010100101011100", "01000110101100001010", "10110110110101001001", "01001110001101010111", "10111010011100101111", "00111010010110100110",
		 "11000010011101101000", "00111110011101010111", "10110110100100001010", "01000110000100001111", "00110010000101011000", "01010110011100110111", "00110110010100100110", "10110010000100111100", "01100110010110101010", "00110010011111010110", "11000010100100010110", "11010010000100111001", "11011110100100111010", "11000110000110000111", "01000010010101101001", "01000110000110001000", "11010010000100110110", "11000011000100111010", "10110010010011111000", "00100011000100100111", "01000110110011111001", "01000110000101111000", "01001010000100101000", "00111010011100001000", "10111010010011110101", "01011010011100000111", "10101110111100100111", "01000001110101010111", "10110110001100000110", "00101101101110011000", "01000010100100110101", "11011010101100011010", "11001110100100011001", "00111001111100011001", "11011001111100100101", "11000010010100111010", "01010010001101001001", "10101010001101011001", "10111011100110010110", "01010010100100000100", "00111110100100100110", "00111101011101000110", "11010001101100100101", "10111101110100111010", "11001110001100111110", "01000101111100010111", "00101101110011000100", "11001001111101110011", "01001010010100010110", "11000010010101000110",
		 "01010010101100101000", "11001001100100100111", "10101110001101001000", "11001010001101111100", "01111010010100111010", "01000010010011111000", "11000010000100011000", "11000101111100000111", "01000010011101110111", "10111111000100101001", "01011010011100110110", "01001101111100100111", "01001010011101010101", "01111010001100001011", "00111110000101010110", "11010010011100111011", "11000010000100011000", "01010101111100001001", "01001010101100000110", "11001110000011100110", "01010110000101010111", "01000010001100001110", "00111010010100100111", "00111010100101011001", "11101010010100010111", "00111001110100111000", "10101010100100011001", "01001110000100010110", "10111010001101000101", "11001101111100010111", "11001110111101000101", "01001010001100011000", "10101101111101011010", "00110010011100010111", "01011110000110100100", "11000110011100011001", "01001110001011101000", "10111001110100111000", "10101101100100011001", "11010110000100010110", "00110011001101000110", "01000011001100100100", "01000101101100001000", "11010011010100000100", "00111110001011010110", "10111110000100110110", "01011110000101000100", "01001010010100101000", "11001110001100011000", "01001110101100010110",
		 "11001110001100001011", "01001010000100100101", "01001110000100101000", "01001010010101000111", "01010001111100110101", "11001010010100000101", "11000110011100010111", "11000110101101011001", "01001110110100010110", "01001111000100000110", "00101001111100011001", "00111010010011001001", "01001101111110010110", "01000110010111001000", "10100110000100011001", "11011110000100011000", "01101101110101010111", "01000110001100110100", "01001010011100011000", "10111110001111001011", "11000010000011111011", "11000010010101100101", "01000010000100010110", "11000110010100010111", "01001010011101110110", "10101001111011101011", "00110110011100111000", "10111101011100100111", "00111010101101000111", "01000010000101011001", "00110010110011011010", "11000010110011101000", "10110001110011110111", "10110110011100110111", "11000110010100001000", "11000010001100110111", "10100101111100001011", "00100010000011101001", "11000110011011101000", "11011111000011100101", "01001010010100100101", "10111010101101011011", "10101010011100110111", "11001110010100001100", "01000010001100100111", "11001110011101111010", "11010010000100010110", "10110010011100011001", "01010001111011100110", "00110110011011000111",
		 "11010010001101001111", "10101010011101001001", "01001110000101001011", "00101010110100111011", "00110001100100000110", "11100111010100010110", "01000110110101111001", "01001010011110001001", "10111101111100100111", "01000110000011001000", "01001101111110011000", "10111010011110101000", "00111110011100001000", "10111010111100101001", "01001101111100010110", "11011111000011101010", "00111111000100111010", "10101010001100110111", "11000011000100001010", "01001110001110010100", "01001001111100110110", "00101110011101110110", "01001010011100110110", "01001001110011100101", "11101010011100111001", "01010110000110001011", "11001110011101111001", "11001001111101000110", "01001111000111000101", "00111010010100000100", "11000010010101111000", "10110110100100010111", "10111110101101110101", "11000111011100101000", "00111110000100001000", "11001110001100101000", "11001011111011111000", "00111010010110010101", "10110110111110010110", "10101110001101000101", "11000010100011101010", "01000010101100111010", "11000010101101111001", "00111110010100010111", "11001010111011110111", "10110010000100000110", "10111010100100011001", "11010110000101101001", "11100101110100111000", "00110010011101000110",
		 "11010010010100110110", "00111010010101011000", "11000010000101010101", "00110001100100000110", "01000110110100010110", "10101010011100000111", "01011010100011001000", "01010110111101001001", "11001010010100101000", "01000010010101101000", "10110110100101001001", "10111010101011110111", "00111110010101011011", "10111110001100100101", "01010010011011101001", "10111001110100000110", "01001010011101010111", "10101110010100110111", "00110110011011100111", "00101001010011111000", "10111110011100101001", "01000010100100000110", "00111010110101001000", "11010110001100110111"); 
				
   data <= weight_ROM(to_integer(unsigned(addr_r)))(to_integer(unsigned(addr_c)));
end arch; 
------------------------------------------------------------------------------------
------ shifter_map1_testbench

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

ENTITY tb_S_MAP1 IS
end tb_S_MAP1;

ARCHITECTURE tb OF tb_S_MAP1 IS

component S_MAP1 is
    GENERIC(
		n : INTEGER := 16;
		addr_col  : integer := 10; -- required bits to store 16 elements
		col : integer := 1023;
        addr_row  : integer := 4; -- required bits to store 16 elements
		row : integer :=12 -- = n
        );
	PORT ( 
		  clk, rst, run: in std_logic;
		  reg_out : out std_logic;
		  din :in std_logic_vector(15 downto 0);
		  df , do , dc ,di : out std_logic_vector (31 downto 0)
		   );
end component;

signal clk, rst, run: std_logic := '1' ;
signal reg_out1 : std_logic ;
signal din1 : std_logic_vector(15 downto 0) := (others => '0');
signal df1 , do1 , dc1 ,di1 : std_logic_vector (31 downto 0);

signal reg_out2 : std_logic ;
signal din2 : std_logic_vector(15 downto 0) := (others => '0');
signal df2 , do2 , dc2 ,di2 : std_logic_vector (31 downto 0);

begin 

map1 : S_MAP1 
    GENERIC MAP(12 , 10 , 1023 , 4 , 12 )
	PORT map( 
		  clk, rst, run,
		  reg_out1,
		  din1 ,
		  df1 , do1 , dc1 ,di1
		   );
		   
map2 : S_MAP1 
    GENERIC MAP(12 , 10 , 1023 , 4 , 12 )
	PORT map( 
		  clk, rst, run,
		  reg_out2,
		  din2 ,
		  df2 , do2 , dc2 ,di2 
		   );
		   
clk <= not clk after 1 ns;
run <= '0' after 10 ns , '1' after 20 ns, '0' after 22 ns;
rst <= '0' after 15 ns;
din1 <= "0101000111101001" after 20 ns, "0111001111101001" after 22 ns, "0101010111101001" after 24 ns, "0101000100101001" after 26 ns, "0101010111001001" after 28 ns, 
	   "0101000101101001" after 30 ns, "0101000110101001" after 32 ns, "0111001100101001" after 34 ns, "0101010110001001" after 36 ns, "0101000110101101" after 38 ns, 
	   "0101010011101001" after 40 ns, "0101100110101001" after 42 ns, "0101010110101001" after 44 ns; 
	   
din2 <= "0100010111101001" after 20 ns, "0011001111101001" after 22 ns, "0001010111101001" after 24 ns, "0100000100101001" after 26 ns, "0001000101101001" after 28 ns, 
	   "0101000111111001" after 30 ns, "0101000011101001" after 32 ns, "0111011111101001" after 34 ns, "0101010111100001" after 36 ns, "0101000100100001" after 38 ns, 
	   "0101010111000001" after 40 ns, "0101000101100001" after 42 ns, "0101000011001001" after 44 ns; 

end tb;
------------------------------------------------------------------------------------
------ shifter_map8_testbench

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

ENTITY tb_S_MAP8 IS
end tb_S_MAP8;

ARCHITECTURE tb OF tb_S_MAP8 IS

component S_MAP1 is
    GENERIC(
		n : INTEGER := 16;
		addr_col  : integer := 10; -- required bits to store 16 elements
		col : integer := 1023;
        addr_row  : integer := 4; -- required bits to store 16 elements
		row : integer :=12 -- = n
        );
	PORT ( 
		  clk, rst, run: in std_logic;
		  reg_out : out std_logic;
		  din :in std_logic_vector(15 downto 0);
		  df , do , dc ,di : out std_logic_vector (31 downto 0)
		   );
end component;

signal clk, rst, run: std_logic := '1' ;
signal din : std_logic_vector(1583 downto 0) := (others => '0');
SIGNAL rego : STD_LOGIC_VECTOR (11 DOWNTO 1 );
SIGNAL data_out_mapf,data_out_mapi,data_out_mapo,data_out_mapg : STD_LOGIC_VECTOR(32*11 -1 DOWNTO 0);

begin 

MAP_1s: FOR I IN 1 TO 11 GENERATE
	MAP1 :  S_MAP1
		GENERIC MAP( 12,
		    10,
		    1023,
			4,
		    12 )
		PORT MAP (  
		    clk,  rst,  run, rego(I),
			din(((I*16)-1) DOWNTO ((I-1)*16)),  
			data_out_mapf((I*32)-1 DOWNTO (I-1)*32),data_out_mapi((I*32)-1 DOWNTO (I-1)*32),
			data_out_mapo((I*32)-1 DOWNTO (I-1)*32),data_out_mapg((I*32)-1 DOWNTO (I-1)*32)
		);
END GENERATE MAP_1s;
		   
clk <= not clk after 1 ns;
--run <= '0' after 10 ns , '1' after 20 ns, '0' after 22 ns ,'1' after  13400 ns, '0' after  13402 ns ;
run <= '0' after 10 ns , '1' after 20 ns, '0' after 22 ns;
rst <= '0' after 15 ns;
--din <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110010101100000101100011110000000000000000000000000000000000000000000000000000000000000000000001101101100000001001101011010000000000000000000001111110001110001001100100101000000000000000000000000000000000000000000000000001101110001010100001100100010000000100111001011000000000000000000001110011111110001010010100010000000000000000000000000000000000000000000000000000100101101001100001100001011000010101110001111000000000000000000001110111101010000010001001010000000000000000000000000000000000000000000000000001110111010101100011000010111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000100000000000000000000000000000000000000000000000000000000000000000011000100001111000000000000000000001110000110100000000000000000000000000000000000000000000000000000000000000000000101101110001100001100011000000000000000000000000000000000000000000000000000000",
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 25 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 27 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000110010110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 29 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111110001000011101100000000000000000000000111100010100000110001011110000000011000010100000000000000000000000000000000000000000000000000000100011001000000101010101010000000000000000000000000000000000000000000000000000001010101011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010010000000100010100000000000000000000000000000000000000000000000000000000000000000000000100000101100000000000000000000000000000000000000000000000000000000000000000000001000111101110100000000000000000000000000000000000000000000000000010000111011010011110111111101000000000000000000011010001110100001000110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 31 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 33 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010110010001010001010100000000000000000000000000000000000000000000000000001001100011010000000000000000000000001111000011000000000000000000000000000000000000000000000000000000000000000000011011101000110000101101100111000000000000000000000000000000000000000000000000000000000000000000001101110010100010000101111110000000000000000000000000000000000000000000000000000011100010110100000000000000000000001011110111000000000000000000010000000000000000000000000000000000000000000000111000101110110000000101110010001001110110111100000000000000000000000000000000000000000000000000110110110110000000011000001010000000000000000000010111100100000000001111100101000000000000000000000000000000000000000000000000" after 35 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011011000011101111100000010110011011010000000000000000000000000000000000001010111011000000001110010101000000000000000000000000000000000000110010011101000110100001111100000000000000000000000000000000000000000000000000001101101100010000100010010000000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 37 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100100110000000000000000000000111101111010000000111100001000000000000000000000000000000000000000000000000000110101110100000001001010101010000111001011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110100111010000000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 39 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 41 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 43 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110111100000000000000000000000000000000000000000000000000000000000000000000000110010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 45 ns,
--	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100110011000000000000000000000000000000000000000000000000000000101011101000000110110111001000000000000000000011100011001000000000000000000000001101101011100000000000000000000000000000000000000000000000000011011101100000000000000000000000000000000000000100110111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101000000000000000000000000000000000000000000000000000000000000000000" after 47 ns;

din <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101111011100010110010110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101001000110001001001100110110001110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100110100001001100101100100000000000000000000000000000000000000000000000000000111100100010000000111001010000000000000000000000000000000000001001011011110000111111100001100000000000000000000000000000000000000000000000000001010011101010000000000000000000000000000000000000000000000000001100101000110000110101010101000010000110000110000000000000000000000000000000000011011010100000001001101111011",
	   "000000000000000000000000000000000001010100100011000100001000100000011110110000100000000000000000000000000000000000000000000000000000000000000000000101011100011100000000000000000001000000110100000001000011101100000000000000000000000000000000000001010000000000111001101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 25 ns,
	   "000000000000000000000000000000000001000010011000001100010110000010100100100001000000000000000000000000000000000000010011001001000000000000000000011000111010110000000000000000000100010100000000011011110000010011000011100001000000000000000000000000000000000001101101011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010000000000000000000000011011111100000000000000000000000000000000000000000000000000000000000000000001100111001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101101011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 27 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101010001110010000001100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000011000011110111010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011011000100110100001000000011101101110000000000000000000000000000000000000000000000000000101001010110000110111101101000000000000000000001000101101110000101100111101000000000000000000000000000000000000000000000000000110100101100100001100110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 29 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101000000000000000000001111111011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000101110000101001000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111100000111100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 31 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 33 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 35 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001000000000000000000000001001110111110000001111100100110000000000000000000000000000000000000000000000000000100100100011000000000000000000010001100001000000000000000000000011100101111000000100101101100000000000000000000000000000000000000101111010010010000101110100000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 37 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010100000000000000000000000000000000000000000000000000000001010010001000000000" after 39 ns,
	   "000000000000010001001101100000000000000000000011010101000000011010111011000000000000000000000000000000000000000000000000000011011110011100000000000000000000000111101010000000000000000000000000000000000000000000000000000000000000000000010001001001001000000000000000000100001001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000110011111010010000001010100111000000000000000000000000000000000000000000000000000001011110100000000000000000000001110000001101000011010110011000000000000000000000000000000000000001001001100100110101001111010000100111110010001011000100111000000000000000000001010100000111000000000000000000000000000000000000000000000000000000000000000000101111101000100000010010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" after 41 ns,
	   "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110010010100000011010000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110001110101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100011110100000100101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011010010000000000000000000000000000000000000000000000000000000000000000000000" after 43 ns,
	   "000000000000000001010110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100100101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011111100000000000000000000000110101011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000101010011011000001010000001000000000000000000000000000000000000000" after 45 ns,
	   "000000000000000010011111001000000000000000000000000101010011000000000000000000000000000000000000001001001000000000000000000000101000000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100111000100000110101010010000000000000000000000000000000000000000000000000000001110011000000000000000000000000001011001111000000000000000000000000000000000000000000000000000000000000000000100001101101110000001000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000010000010010000101010000101101101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010111110000000010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100100000000000000000000000000000000000000000000000000000000000000000000" after 47 ns;

PROCESS
BEGIN
	REPORT " The first outputs are :\n out_f = " & integer'image(to_integer(signed(data_out_mapf))) & "\n out_i = " & integer'image(to_integer(signed(data_out_mapi))) &  
		   ":\n out_o = " & integer'image(to_integer(signed(data_out_mapo))) & "\n out_g = " & integer'image(to_integer(signed(data_out_mapg)))
		   SEVERITY NOTE;
	WAIT FOR 370 NS;
	WAIT;
END PROCESS;

--din <= "",
--	   "" after 25 ns,
--	   "" after 27 ns,
--	   "" after 29 ns,
--	   "" after 31 ns,
--	   "" after 33 ns,
--	   "" after 35 ns,
--	   "" after 37 ns,
--	   "" after 39 ns,
--	   "" after 41 ns,
--	   "" after 43 ns,
--	   "" after 45 ns,
--	   "" after 47 ns;
end tb;
